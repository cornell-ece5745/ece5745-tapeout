magic
tech sky130A
magscale 1 2
timestamp 1655409329
<< obsli1 >>
rect 1104 2159 178848 177361
<< obsm1 >>
rect 14 2128 179754 177392
<< metal2 >>
rect 23846 179200 23902 180000
rect 63130 179200 63186 180000
rect 101770 179200 101826 180000
rect 141054 179200 141110 180000
rect 179694 179200 179750 180000
rect 18 0 74 800
rect 38658 0 38714 800
rect 77942 0 77998 800
rect 116582 0 116638 800
rect 155866 0 155922 800
<< obsm2 >>
rect 20 179144 23790 179330
rect 23958 179144 63074 179330
rect 63242 179144 101714 179330
rect 101882 179144 140998 179330
rect 141166 179144 179638 179330
rect 20 856 179748 179144
rect 130 800 38602 856
rect 38770 800 77886 856
rect 78054 800 116526 856
rect 116694 800 155810 856
rect 155978 800 179748 856
<< metal3 >>
rect 0 164568 800 164688
rect 179200 138728 180000 138848
rect 0 123088 800 123208
rect 179200 97248 180000 97368
rect 0 82288 800 82408
rect 179200 56448 180000 56568
rect 0 40808 800 40928
rect 179200 14968 180000 15088
<< obsm3 >>
rect 800 164768 179200 177377
rect 880 164488 179200 164768
rect 800 138928 179200 164488
rect 800 138648 179120 138928
rect 800 123288 179200 138648
rect 880 123008 179200 123288
rect 800 97448 179200 123008
rect 800 97168 179120 97448
rect 800 82488 179200 97168
rect 880 82208 179200 82488
rect 800 56648 179200 82208
rect 800 56368 179120 56648
rect 800 41008 179200 56368
rect 880 40728 179200 41008
rect 800 15168 179200 40728
rect 800 14888 179120 15168
rect 800 2143 179200 14888
<< metal4 >>
rect 4208 2128 4528 177392
rect 19568 2128 19888 177392
rect 34928 2128 35248 177392
rect 50288 2128 50608 177392
rect 65648 2128 65968 177392
rect 81008 2128 81328 177392
rect 96368 2128 96688 177392
rect 111728 2128 112048 177392
rect 127088 2128 127408 177392
rect 142448 2128 142768 177392
rect 157808 2128 158128 177392
rect 173168 2128 173488 177392
<< obsm4 >>
rect 67403 70891 80928 129845
rect 81408 70891 96288 129845
rect 96768 70891 111648 129845
rect 112128 70891 127008 129845
rect 127488 70891 136101 129845
<< labels >>
rlabel metal3 s 179200 14968 180000 15088 6 adapter_parity
port 1 nsew signal output
rlabel metal3 s 179200 138728 180000 138848 6 ap_en
port 2 nsew signal output
rlabel metal2 s 101770 179200 101826 180000 6 clk
port 3 nsew signal input
rlabel metal2 s 116582 0 116638 800 6 clk_en
port 4 nsew signal output
rlabel metal3 s 0 164568 800 164688 6 cs_en
port 5 nsew signal output
rlabel metal2 s 63130 179200 63186 180000 6 loopthrough_sel
port 6 nsew signal input
rlabel metal2 s 18 0 74 800 6 lt_sel_en
port 7 nsew signal output
rlabel metal2 s 179694 179200 179750 180000 6 minion_parity
port 8 nsew signal output
rlabel metal2 s 155866 0 155922 800 6 miso_en
port 9 nsew signal output
rlabel metal2 s 38658 0 38714 800 6 mosi_en
port 10 nsew signal output
rlabel metal3 s 0 40808 800 40928 6 mp_en
port 11 nsew signal output
rlabel metal3 s 179200 97248 180000 97368 6 reset
port 12 nsew signal input
rlabel metal3 s 0 82288 800 82408 6 reset_en
port 13 nsew signal output
rlabel metal2 s 141054 179200 141110 180000 6 sclk_en
port 14 nsew signal output
rlabel metal2 s 77942 0 77998 800 6 spi_min_cs
port 15 nsew signal input
rlabel metal3 s 0 123088 800 123208 6 spi_min_miso
port 16 nsew signal output
rlabel metal2 s 23846 179200 23902 180000 6 spi_min_mosi
port 17 nsew signal input
rlabel metal3 s 179200 56448 180000 56568 6 spi_min_sclk
port 18 nsew signal input
rlabel metal4 s 4208 2128 4528 177392 6 vccd1
port 19 nsew power input
rlabel metal4 s 34928 2128 35248 177392 6 vccd1
port 19 nsew power input
rlabel metal4 s 65648 2128 65968 177392 6 vccd1
port 19 nsew power input
rlabel metal4 s 96368 2128 96688 177392 6 vccd1
port 19 nsew power input
rlabel metal4 s 127088 2128 127408 177392 6 vccd1
port 19 nsew power input
rlabel metal4 s 157808 2128 158128 177392 6 vccd1
port 19 nsew power input
rlabel metal4 s 19568 2128 19888 177392 6 vssd1
port 20 nsew ground input
rlabel metal4 s 50288 2128 50608 177392 6 vssd1
port 20 nsew ground input
rlabel metal4 s 81008 2128 81328 177392 6 vssd1
port 20 nsew ground input
rlabel metal4 s 111728 2128 112048 177392 6 vssd1
port 20 nsew ground input
rlabel metal4 s 142448 2128 142768 177392 6 vssd1
port 20 nsew ground input
rlabel metal4 s 173168 2128 173488 177392 6 vssd1
port 20 nsew ground input
<< properties >>
string FIXED_BBOX 0 0 180000 180000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 18895134
string GDS_FILE /home/acm289/ece5745-tapeout/openlane/project-group15/runs/project-group15/results/finishing/grp_15_SPI_TapeOutBlockRTL_32bits_5entries.magic.gds
string GDS_START 625260
<< end >>


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO grp_99_SPI_TapeOutBlockRTL_32bits_5entries
  CLASS BLOCK ;
  FOREIGN grp_99_SPI_TapeOutBlockRTL_32bits_5entries ;
  ORIGIN 0.000 0.000 ;
  SIZE 1210.000 BY 1510.000 ;
  PIN adapter_parity
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 604.990 1506.000 605.270 1510.000 ;
    END
  END adapter_parity
  PIN ap_en
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 777.030 0.000 777.310 4.000 ;
    END
  END ap_en
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.110 0.000 86.390 4.000 ;
    END
  END clk
  PIN clk_en
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 258.610 0.000 258.890 4.000 ;
    END
  END clk_en
  PIN cs_en
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1206.000 188.400 1210.000 189.000 ;
    END
  END cs_en
  PIN loopthrough_sel
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.070 1506.000 121.350 1510.000 ;
    END
  END loopthrough_sel
  PIN lt_sel_en
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 846.950 1506.000 847.230 1510.000 ;
    END
  END lt_sel_en
  PIN minion_parity
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.030 1506.000 363.310 1510.000 ;
    END
  END minion_parity
  PIN miso_en
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1206.000 565.800 1210.000 566.400 ;
    END
  END miso_en
  PIN mosi_en
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1206.000 943.200 1210.000 943.800 ;
    END
  END mosi_en
  PIN mp_en
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 377.440 4.000 378.040 ;
    END
  END mp_en
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 431.570 0.000 431.850 4.000 ;
    END
  END reset
  PIN reset_en
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 604.530 0.000 604.810 4.000 ;
    END
  END reset_en
  PIN sclk_en
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1206.000 1320.600 1210.000 1321.200 ;
    END
  END sclk_en
  PIN spi_min__cs
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1088.910 1506.000 1089.190 1510.000 ;
    END
  END spi_min__cs
  PIN spi_min__miso
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 949.990 0.000 950.270 4.000 ;
    END
  END spi_min__miso
  PIN spi_min__mosi
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1132.240 4.000 1132.840 ;
    END
  END spi_min__mosi
  PIN spi_min__sclk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1122.950 0.000 1123.230 4.000 ;
    END
  END spi_min__sclk
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 1498.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 1498.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 1498.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 1498.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 1498.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 1498.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 942.640 10.640 944.240 1498.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 1096.240 10.640 1097.840 1498.960 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 1498.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 1498.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 1498.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 1498.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 1498.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 1498.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 1019.440 10.640 1021.040 1498.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 1173.040 10.640 1174.640 1498.960 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 1204.280 1498.805 ;
      LAYER met1 ;
        RECT 5.520 10.640 1204.280 1498.960 ;
      LAYER met2 ;
        RECT 6.990 1505.720 120.790 1506.610 ;
        RECT 121.630 1505.720 362.750 1506.610 ;
        RECT 363.590 1505.720 604.710 1506.610 ;
        RECT 605.550 1505.720 846.670 1506.610 ;
        RECT 847.510 1505.720 1088.630 1506.610 ;
        RECT 1089.470 1505.720 1200.970 1506.610 ;
        RECT 6.990 4.280 1200.970 1505.720 ;
        RECT 6.990 4.000 85.830 4.280 ;
        RECT 86.670 4.000 258.330 4.280 ;
        RECT 259.170 4.000 431.290 4.280 ;
        RECT 432.130 4.000 604.250 4.280 ;
        RECT 605.090 4.000 776.750 4.280 ;
        RECT 777.590 4.000 949.710 4.280 ;
        RECT 950.550 4.000 1122.670 4.280 ;
        RECT 1123.510 4.000 1200.970 4.280 ;
      LAYER met3 ;
        RECT 4.000 1321.600 1206.000 1498.885 ;
        RECT 4.000 1320.200 1205.600 1321.600 ;
        RECT 4.000 1133.240 1206.000 1320.200 ;
        RECT 4.400 1131.840 1206.000 1133.240 ;
        RECT 4.000 944.200 1206.000 1131.840 ;
        RECT 4.000 942.800 1205.600 944.200 ;
        RECT 4.000 566.800 1206.000 942.800 ;
        RECT 4.000 565.400 1205.600 566.800 ;
        RECT 4.000 378.440 1206.000 565.400 ;
        RECT 4.400 377.040 1206.000 378.440 ;
        RECT 4.000 189.400 1206.000 377.040 ;
        RECT 4.000 188.000 1205.600 189.400 ;
        RECT 4.000 10.715 1206.000 188.000 ;
      LAYER met4 ;
        RECT 484.215 673.375 558.240 1001.465 ;
        RECT 560.640 673.375 635.040 1001.465 ;
        RECT 637.440 673.375 711.840 1001.465 ;
        RECT 714.240 673.375 778.945 1001.465 ;
  END
END grp_99_SPI_TapeOutBlockRTL_32bits_5entries
END LIBRARY


magic
tech sky130A
magscale 1 2
timestamp 1654617189
<< obsli1 >>
rect 1104 2159 240856 299761
<< obsm1 >>
rect 1104 2128 240856 299792
<< metal2 >>
rect 40314 301200 40370 302000
rect 120906 301200 120962 302000
rect 201590 301200 201646 302000
rect 17222 0 17278 800
rect 51722 0 51778 800
rect 86314 0 86370 800
rect 120906 0 120962 800
rect 155406 0 155462 800
rect 189998 0 190054 800
rect 224590 0 224646 800
<< obsm2 >>
rect 1398 301144 40258 301322
rect 40426 301144 120850 301322
rect 121018 301144 201534 301322
rect 201702 301144 240194 301322
rect 1398 856 240194 301144
rect 1398 734 17166 856
rect 17334 734 51666 856
rect 51834 734 86258 856
rect 86426 734 120850 856
rect 121018 734 155350 856
rect 155518 734 189942 856
rect 190110 734 224534 856
rect 224702 734 240194 856
<< metal3 >>
rect 241200 280304 242000 280424
rect 241200 237192 242000 237312
rect 241200 194080 242000 194200
rect 0 150968 800 151088
rect 241200 150832 242000 150952
rect 241200 107720 242000 107840
rect 241200 64608 242000 64728
rect 241200 21496 242000 21616
<< obsm3 >>
rect 800 280504 241200 299777
rect 800 280224 241120 280504
rect 800 237392 241200 280224
rect 800 237112 241120 237392
rect 800 194280 241200 237112
rect 800 194000 241120 194280
rect 800 151168 241200 194000
rect 880 151032 241200 151168
rect 880 150888 241120 151032
rect 800 150752 241120 150888
rect 800 107920 241200 150752
rect 800 107640 241120 107920
rect 800 64808 241200 107640
rect 800 64528 241120 64808
rect 800 21696 241200 64528
rect 800 21416 241120 21696
rect 800 2143 241200 21416
<< metal4 >>
rect 4208 2128 4528 299792
rect 19568 2128 19888 299792
rect 34928 2128 35248 299792
rect 50288 2128 50608 299792
rect 65648 2128 65968 299792
rect 81008 2128 81328 299792
rect 96368 2128 96688 299792
rect 111728 2128 112048 299792
rect 127088 2128 127408 299792
rect 142448 2128 142768 299792
rect 157808 2128 158128 299792
rect 173168 2128 173488 299792
rect 188528 2128 188848 299792
rect 203888 2128 204208 299792
rect 219248 2128 219568 299792
rect 234608 2128 234928 299792
<< obsm4 >>
rect 133643 126379 142368 189141
rect 142848 126379 157728 189141
rect 158208 126379 173088 189141
rect 173568 126379 188448 189141
rect 188928 126379 203808 189141
rect 204288 126379 209333 189141
<< labels >>
rlabel metal2 s 201590 301200 201646 302000 6 adapter_parity
port 1 nsew signal output
rlabel metal3 s 241200 194080 242000 194200 6 ap_en
port 2 nsew signal output
rlabel metal2 s 17222 0 17278 800 6 clk
port 3 nsew signal input
rlabel metal2 s 51722 0 51778 800 6 clk_en
port 4 nsew signal output
rlabel metal3 s 241200 21496 242000 21616 6 cs_en
port 5 nsew signal output
rlabel metal2 s 40314 301200 40370 302000 6 loopthrough_sel
port 6 nsew signal input
rlabel metal3 s 0 150968 800 151088 6 lt_sel_en
port 7 nsew signal output
rlabel metal2 s 120906 301200 120962 302000 6 minion_parity
port 8 nsew signal output
rlabel metal3 s 241200 64608 242000 64728 6 miso_en
port 9 nsew signal output
rlabel metal3 s 241200 107720 242000 107840 6 mosi_en
port 10 nsew signal output
rlabel metal3 s 241200 237192 242000 237312 6 mp_en
port 11 nsew signal output
rlabel metal2 s 86314 0 86370 800 6 reset
port 12 nsew signal input
rlabel metal2 s 120906 0 120962 800 6 reset_en
port 13 nsew signal output
rlabel metal3 s 241200 150832 242000 150952 6 sclk_en
port 14 nsew signal output
rlabel metal2 s 155406 0 155462 800 6 spi_min__cs
port 15 nsew signal input
rlabel metal3 s 241200 280304 242000 280424 6 spi_min__miso
port 16 nsew signal output
rlabel metal2 s 189998 0 190054 800 6 spi_min__mosi
port 17 nsew signal input
rlabel metal2 s 224590 0 224646 800 6 spi_min__sclk
port 18 nsew signal input
rlabel metal4 s 4208 2128 4528 299792 6 vccd1
port 19 nsew power input
rlabel metal4 s 34928 2128 35248 299792 6 vccd1
port 19 nsew power input
rlabel metal4 s 65648 2128 65968 299792 6 vccd1
port 19 nsew power input
rlabel metal4 s 96368 2128 96688 299792 6 vccd1
port 19 nsew power input
rlabel metal4 s 127088 2128 127408 299792 6 vccd1
port 19 nsew power input
rlabel metal4 s 157808 2128 158128 299792 6 vccd1
port 19 nsew power input
rlabel metal4 s 188528 2128 188848 299792 6 vccd1
port 19 nsew power input
rlabel metal4 s 219248 2128 219568 299792 6 vccd1
port 19 nsew power input
rlabel metal4 s 19568 2128 19888 299792 6 vssd1
port 20 nsew ground input
rlabel metal4 s 50288 2128 50608 299792 6 vssd1
port 20 nsew ground input
rlabel metal4 s 81008 2128 81328 299792 6 vssd1
port 20 nsew ground input
rlabel metal4 s 111728 2128 112048 299792 6 vssd1
port 20 nsew ground input
rlabel metal4 s 142448 2128 142768 299792 6 vssd1
port 20 nsew ground input
rlabel metal4 s 173168 2128 173488 299792 6 vssd1
port 20 nsew ground input
rlabel metal4 s 203888 2128 204208 299792 6 vssd1
port 20 nsew ground input
rlabel metal4 s 234608 2128 234928 299792 6 vssd1
port 20 nsew ground input
<< properties >>
string FIXED_BBOX 0 0 242000 302000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 28443730
string GDS_FILE /home/acm289/ece5745-tapeout/openlane/project-group99/runs/project-group99/results/finishing/grp_99_SPI_TapeOutBlockRTL_32bits_5entries.magic.gds
string GDS_START 487654
<< end >>


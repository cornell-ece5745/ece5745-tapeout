magic
tech sky130A
magscale 1 2
timestamp 1655334262
<< obsli1 >>
rect 1104 2159 240856 299761
<< obsm1 >>
rect 1104 2128 240856 299792
<< metal2 >>
rect 20166 301200 20222 302000
rect 60462 301200 60518 302000
rect 100758 301200 100814 302000
rect 141146 301200 141202 302000
rect 181442 301200 181498 302000
rect 221738 301200 221794 302000
rect 30194 0 30250 800
rect 90638 0 90694 800
rect 151174 0 151230 800
rect 211618 0 211674 800
<< obsm2 >>
rect 1398 301144 20110 301322
rect 20278 301144 60406 301322
rect 60574 301144 100702 301322
rect 100870 301144 141090 301322
rect 141258 301144 181386 301322
rect 181554 301144 221682 301322
rect 221850 301144 240194 301322
rect 1398 856 240194 301144
rect 1398 734 30138 856
rect 30306 734 90582 856
rect 90750 734 151118 856
rect 151286 734 211562 856
rect 211730 734 240194 856
<< metal3 >>
rect 241200 280304 242000 280424
rect 241200 237192 242000 237312
rect 241200 194080 242000 194200
rect 0 150968 800 151088
rect 241200 150832 242000 150952
rect 241200 107720 242000 107840
rect 241200 64608 242000 64728
rect 241200 21496 242000 21616
<< obsm3 >>
rect 800 280504 241200 299777
rect 800 280224 241120 280504
rect 800 237392 241200 280224
rect 800 237112 241120 237392
rect 800 194280 241200 237112
rect 800 194000 241120 194280
rect 800 151168 241200 194000
rect 880 151032 241200 151168
rect 880 150888 241120 151032
rect 800 150752 241120 150888
rect 800 107920 241200 150752
rect 800 107640 241120 107920
rect 800 64808 241200 107640
rect 800 64528 241120 64808
rect 800 21696 241200 64528
rect 800 21416 241120 21696
rect 800 2143 241200 21416
<< metal4 >>
rect 4208 2128 4528 299792
rect 19568 2128 19888 299792
rect 34928 2128 35248 299792
rect 50288 2128 50608 299792
rect 65648 2128 65968 299792
rect 81008 2128 81328 299792
rect 96368 2128 96688 299792
rect 111728 2128 112048 299792
rect 127088 2128 127408 299792
rect 142448 2128 142768 299792
rect 157808 2128 158128 299792
rect 173168 2128 173488 299792
rect 188528 2128 188848 299792
rect 203888 2128 204208 299792
rect 219248 2128 219568 299792
rect 234608 2128 234928 299792
<< obsm4 >>
rect 97763 212331 111648 276997
rect 112128 212331 127008 276997
rect 127488 212331 142368 276997
rect 142848 212331 157728 276997
rect 158208 212331 173088 276997
rect 173568 212331 174557 276997
<< labels >>
rlabel metal2 s 100758 301200 100814 302000 6 adapter_parity
port 1 nsew signal output
rlabel metal3 s 0 150968 800 151088 6 ap_en
port 2 nsew signal output
rlabel metal2 s 30194 0 30250 800 6 clk
port 3 nsew signal input
rlabel metal2 s 90638 0 90694 800 6 clk_en
port 4 nsew signal output
rlabel metal3 s 241200 21496 242000 21616 6 cs_en
port 5 nsew signal output
rlabel metal2 s 20166 301200 20222 302000 6 loopthrough_sel
port 6 nsew signal input
rlabel metal3 s 241200 194080 242000 194200 6 lt_sel_en
port 7 nsew signal output
rlabel metal2 s 60462 301200 60518 302000 6 minion_parity
port 8 nsew signal output
rlabel metal3 s 241200 64608 242000 64728 6 miso_en
port 9 nsew signal output
rlabel metal3 s 241200 107720 242000 107840 6 mosi_en
port 10 nsew signal output
rlabel metal2 s 141146 301200 141202 302000 6 mp_en
port 11 nsew signal output
rlabel metal2 s 151174 0 151230 800 6 reset
port 12 nsew signal input
rlabel metal2 s 211618 0 211674 800 6 reset_en
port 13 nsew signal output
rlabel metal3 s 241200 150832 242000 150952 6 sclk_en
port 14 nsew signal output
rlabel metal2 s 181442 301200 181498 302000 6 spi_min_cs
port 15 nsew signal input
rlabel metal3 s 241200 237192 242000 237312 6 spi_min_miso
port 16 nsew signal output
rlabel metal3 s 241200 280304 242000 280424 6 spi_min_mosi
port 17 nsew signal input
rlabel metal2 s 221738 301200 221794 302000 6 spi_min_sclk
port 18 nsew signal input
rlabel metal4 s 4208 2128 4528 299792 6 vccd1
port 19 nsew power input
rlabel metal4 s 34928 2128 35248 299792 6 vccd1
port 19 nsew power input
rlabel metal4 s 65648 2128 65968 299792 6 vccd1
port 19 nsew power input
rlabel metal4 s 96368 2128 96688 299792 6 vccd1
port 19 nsew power input
rlabel metal4 s 127088 2128 127408 299792 6 vccd1
port 19 nsew power input
rlabel metal4 s 157808 2128 158128 299792 6 vccd1
port 19 nsew power input
rlabel metal4 s 188528 2128 188848 299792 6 vccd1
port 19 nsew power input
rlabel metal4 s 219248 2128 219568 299792 6 vccd1
port 19 nsew power input
rlabel metal4 s 19568 2128 19888 299792 6 vssd1
port 20 nsew ground input
rlabel metal4 s 50288 2128 50608 299792 6 vssd1
port 20 nsew ground input
rlabel metal4 s 81008 2128 81328 299792 6 vssd1
port 20 nsew ground input
rlabel metal4 s 111728 2128 112048 299792 6 vssd1
port 20 nsew ground input
rlabel metal4 s 142448 2128 142768 299792 6 vssd1
port 20 nsew ground input
rlabel metal4 s 173168 2128 173488 299792 6 vssd1
port 20 nsew ground input
rlabel metal4 s 203888 2128 204208 299792 6 vssd1
port 20 nsew ground input
rlabel metal4 s 234608 2128 234928 299792 6 vssd1
port 20 nsew ground input
<< properties >>
string FIXED_BBOX 0 0 242000 302000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 29642224
string GDS_FILE /home/acm289/ece5745-tapeout/openlane/project-group99/runs/project-group99/results/finishing/grp_99_SPI_TapeOutBlockRTL_32bits_5entries.magic.gds
string GDS_START 599388
<< end >>


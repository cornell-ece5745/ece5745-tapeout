magic
tech sky130A
magscale 1 2
timestamp 1655489412
<< obsli1 >>
rect 1104 2159 138828 137649
<< obsm1 >>
rect 1104 2128 138828 137680
<< metal2 >>
rect 11610 139200 11666 140000
rect 34886 139200 34942 140000
rect 58254 139200 58310 140000
rect 81622 139200 81678 140000
rect 104898 139200 104954 140000
rect 128266 139200 128322 140000
rect 9954 0 10010 800
rect 29918 0 29974 800
rect 49882 0 49938 800
rect 69938 0 69994 800
rect 89902 0 89958 800
rect 109958 0 110014 800
rect 129922 0 129978 800
<< obsm2 >>
rect 1398 139144 11554 139346
rect 11722 139144 34830 139346
rect 34998 139144 58198 139346
rect 58366 139144 81566 139346
rect 81734 139144 104842 139346
rect 105010 139144 128210 139346
rect 128378 139144 138164 139346
rect 1398 856 138164 139144
rect 1398 800 9898 856
rect 10066 800 29862 856
rect 30030 800 49826 856
rect 49994 800 69882 856
rect 70050 800 89846 856
rect 90014 800 109902 856
rect 110070 800 129866 856
rect 130034 800 138164 856
<< metal3 >>
rect 0 125808 800 125928
rect 0 97792 800 97912
rect 0 69776 800 69896
rect 0 41760 800 41880
rect 0 13880 800 14000
<< obsm3 >>
rect 800 126008 136699 137665
rect 880 125728 136699 126008
rect 800 97992 136699 125728
rect 880 97712 136699 97992
rect 800 69976 136699 97712
rect 880 69696 136699 69976
rect 800 41960 136699 69696
rect 880 41680 136699 41960
rect 800 14080 136699 41680
rect 880 13800 136699 14080
rect 800 2143 136699 13800
<< metal4 >>
rect 4208 2128 4528 137680
rect 19568 2128 19888 137680
rect 34928 2128 35248 137680
rect 50288 2128 50608 137680
rect 65648 2128 65968 137680
rect 81008 2128 81328 137680
rect 96368 2128 96688 137680
rect 111728 2128 112048 137680
rect 127088 2128 127408 137680
<< obsm4 >>
rect 22691 2483 34848 126309
rect 35328 2483 50208 126309
rect 50688 2483 65568 126309
rect 66048 2483 80928 126309
rect 81408 2483 96288 126309
rect 96768 2483 111648 126309
rect 112128 2483 126901 126309
<< labels >>
rlabel metal2 s 49882 0 49938 800 6 adapter_parity
port 1 nsew signal output
rlabel metal2 s 69938 0 69994 800 6 ap_en
port 2 nsew signal output
rlabel metal2 s 11610 139200 11666 140000 6 clk
port 3 nsew signal input
rlabel metal2 s 34886 139200 34942 140000 6 clk_en
port 4 nsew signal output
rlabel metal2 s 104898 139200 104954 140000 6 cs_en
port 5 nsew signal output
rlabel metal3 s 0 69776 800 69896 6 loopthrough_sel
port 6 nsew signal input
rlabel metal2 s 89902 0 89958 800 6 lt_sel_en
port 7 nsew signal output
rlabel metal3 s 0 97792 800 97912 6 minion_parity
port 8 nsew signal output
rlabel metal2 s 128266 139200 128322 140000 6 miso_en
port 9 nsew signal output
rlabel metal3 s 0 125808 800 125928 6 mosi_en
port 10 nsew signal output
rlabel metal2 s 109958 0 110014 800 6 mp_en
port 11 nsew signal output
rlabel metal2 s 58254 139200 58310 140000 6 reset
port 12 nsew signal input
rlabel metal2 s 81622 139200 81678 140000 6 reset_en
port 13 nsew signal output
rlabel metal2 s 129922 0 129978 800 6 sclk_en
port 14 nsew signal output
rlabel metal2 s 29918 0 29974 800 6 spi_min_cs
port 15 nsew signal input
rlabel metal3 s 0 13880 800 14000 6 spi_min_miso
port 16 nsew signal output
rlabel metal3 s 0 41760 800 41880 6 spi_min_mosi
port 17 nsew signal input
rlabel metal2 s 9954 0 10010 800 6 spi_min_sclk
port 18 nsew signal input
rlabel metal4 s 4208 2128 4528 137680 6 vccd1
port 19 nsew power input
rlabel metal4 s 34928 2128 35248 137680 6 vccd1
port 19 nsew power input
rlabel metal4 s 65648 2128 65968 137680 6 vccd1
port 19 nsew power input
rlabel metal4 s 96368 2128 96688 137680 6 vccd1
port 19 nsew power input
rlabel metal4 s 127088 2128 127408 137680 6 vccd1
port 19 nsew power input
rlabel metal4 s 19568 2128 19888 137680 6 vssd1
port 20 nsew ground input
rlabel metal4 s 50288 2128 50608 137680 6 vssd1
port 20 nsew ground input
rlabel metal4 s 81008 2128 81328 137680 6 vssd1
port 20 nsew ground input
rlabel metal4 s 111728 2128 112048 137680 6 vssd1
port 20 nsew ground input
<< properties >>
string FIXED_BBOX 0 0 140000 140000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 31334106
string GDS_FILE /home/acm289/ece5745-tapeout/openlane/project-group17/runs/project-group17/results/finishing/grp_17_SPI_TapeOutBlockRTL_32bits_5entries.magic.gds
string GDS_START 1333880
<< end >>


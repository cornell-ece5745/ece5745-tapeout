VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO grp_99_SPI_TapeOutBlockRTL_32bits_5entries
  CLASS BLOCK ;
  FOREIGN grp_99_SPI_TapeOutBlockRTL_32bits_5entries ;
  ORIGIN 0.000 0.000 ;
  SIZE 1210.000 BY 1510.000 ;
  PIN adapter_parity
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1007.950 1506.000 1008.230 1510.000 ;
    END
  END adapter_parity
  PIN ap_en
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 907.210 0.000 907.490 4.000 ;
    END
  END ap_en
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 100.830 0.000 101.110 4.000 ;
    END
  END clk
  PIN clk_en
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 302.310 0.000 302.590 4.000 ;
    END
  END clk_en
  PIN cs_en
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1206.000 125.840 1210.000 126.440 ;
    END
  END cs_en
  PIN loopthrough_sel
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 201.570 1506.000 201.850 1510.000 ;
    END
  END loopthrough_sel
  PIN lt_sel_en
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 251.640 4.000 252.240 ;
    END
  END lt_sel_en
  PIN minion_parity
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 604.530 1506.000 604.810 1510.000 ;
    END
  END minion_parity
  PIN miso_en
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1206.000 377.440 1210.000 378.040 ;
    END
  END miso_en
  PIN mosi_en
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1206.000 629.040 1210.000 629.640 ;
    END
  END mosi_en
  PIN mp_en
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 754.840 4.000 755.440 ;
    END
  END mp_en
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 503.790 0.000 504.070 4.000 ;
    END
  END reset
  PIN reset_en
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 705.730 0.000 706.010 4.000 ;
    END
  END reset_en
  PIN sclk_en
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1206.000 880.640 1210.000 881.240 ;
    END
  END sclk_en
  PIN spi_min__cs
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1206.000 1132.240 1210.000 1132.840 ;
    END
  END spi_min__cs
  PIN spi_min__miso
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1108.690 0.000 1108.970 4.000 ;
    END
  END spi_min__miso
  PIN spi_min__mosi
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1258.040 4.000 1258.640 ;
    END
  END spi_min__mosi
  PIN spi_min__sclk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1206.000 1383.840 1210.000 1384.440 ;
    END
  END spi_min__sclk
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 1498.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 1498.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 1498.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 1498.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 1498.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 1498.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 942.640 10.640 944.240 1498.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 1096.240 10.640 1097.840 1498.960 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 1498.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 1498.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 1498.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 1498.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 1498.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 1498.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 1019.440 10.640 1021.040 1498.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 1173.040 10.640 1174.640 1498.960 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 1204.280 1498.805 ;
      LAYER met1 ;
        RECT 5.520 10.640 1204.280 1498.960 ;
      LAYER met2 ;
        RECT 6.990 1505.720 201.290 1506.610 ;
        RECT 202.130 1505.720 604.250 1506.610 ;
        RECT 605.090 1505.720 1007.670 1506.610 ;
        RECT 1008.510 1505.720 1200.970 1506.610 ;
        RECT 6.990 4.280 1200.970 1505.720 ;
        RECT 6.990 3.670 100.550 4.280 ;
        RECT 101.390 3.670 302.030 4.280 ;
        RECT 302.870 3.670 503.510 4.280 ;
        RECT 504.350 3.670 705.450 4.280 ;
        RECT 706.290 3.670 906.930 4.280 ;
        RECT 907.770 3.670 1108.410 4.280 ;
        RECT 1109.250 3.670 1200.970 4.280 ;
      LAYER met3 ;
        RECT 4.000 1384.840 1206.000 1498.885 ;
        RECT 4.000 1383.440 1205.600 1384.840 ;
        RECT 4.000 1259.040 1206.000 1383.440 ;
        RECT 4.400 1257.640 1206.000 1259.040 ;
        RECT 4.000 1133.240 1206.000 1257.640 ;
        RECT 4.000 1131.840 1205.600 1133.240 ;
        RECT 4.000 881.640 1206.000 1131.840 ;
        RECT 4.000 880.240 1205.600 881.640 ;
        RECT 4.000 755.840 1206.000 880.240 ;
        RECT 4.400 754.440 1206.000 755.840 ;
        RECT 4.000 630.040 1206.000 754.440 ;
        RECT 4.000 628.640 1205.600 630.040 ;
        RECT 4.000 378.440 1206.000 628.640 ;
        RECT 4.000 377.040 1205.600 378.440 ;
        RECT 4.000 252.640 1206.000 377.040 ;
        RECT 4.400 251.240 1206.000 252.640 ;
        RECT 4.000 126.840 1206.000 251.240 ;
        RECT 4.000 125.440 1205.600 126.840 ;
        RECT 4.000 10.715 1206.000 125.440 ;
      LAYER met4 ;
        RECT 510.895 703.295 558.240 1168.745 ;
        RECT 560.640 703.295 635.040 1168.745 ;
        RECT 637.440 703.295 711.840 1168.745 ;
        RECT 714.240 703.295 788.640 1168.745 ;
        RECT 791.040 703.295 865.440 1168.745 ;
        RECT 867.840 703.295 879.225 1168.745 ;
  END
END grp_99_SPI_TapeOutBlockRTL_32bits_5entries
END LIBRARY


magic
tech sky130A
magscale 1 2
timestamp 1654995097
<< obsli1 >>
rect 1104 2159 240856 299761
<< obsm1 >>
rect 1104 2128 240856 299792
<< metal2 >>
rect 24214 301200 24270 302000
rect 72606 301200 72662 302000
rect 120998 301200 121054 302000
rect 169390 301200 169446 302000
rect 217782 301200 217838 302000
rect 17222 0 17278 800
rect 51722 0 51778 800
rect 86314 0 86370 800
rect 120906 0 120962 800
rect 155406 0 155462 800
rect 189998 0 190054 800
rect 224590 0 224646 800
<< obsm2 >>
rect 1398 301144 24158 301322
rect 24326 301144 72550 301322
rect 72718 301144 120942 301322
rect 121110 301144 169334 301322
rect 169502 301144 217726 301322
rect 217894 301144 240194 301322
rect 1398 856 240194 301144
rect 1398 800 17166 856
rect 17334 800 51666 856
rect 51834 800 86258 856
rect 86426 800 120850 856
rect 121018 800 155350 856
rect 155518 800 189942 856
rect 190110 800 224534 856
rect 224702 800 240194 856
<< metal3 >>
rect 241200 264120 242000 264240
rect 0 226448 800 226568
rect 241200 188640 242000 188760
rect 241200 113160 242000 113280
rect 0 75488 800 75608
rect 241200 37680 242000 37800
<< obsm3 >>
rect 800 264320 241200 299777
rect 800 264040 241120 264320
rect 800 226648 241200 264040
rect 880 226368 241200 226648
rect 800 188840 241200 226368
rect 800 188560 241120 188840
rect 800 113360 241200 188560
rect 800 113080 241120 113360
rect 800 75688 241200 113080
rect 880 75408 241200 75688
rect 800 37880 241200 75408
rect 800 37600 241120 37880
rect 800 2143 241200 37600
<< metal4 >>
rect 4208 2128 4528 299792
rect 19568 2128 19888 299792
rect 34928 2128 35248 299792
rect 50288 2128 50608 299792
rect 65648 2128 65968 299792
rect 81008 2128 81328 299792
rect 96368 2128 96688 299792
rect 111728 2128 112048 299792
rect 127088 2128 127408 299792
rect 142448 2128 142768 299792
rect 157808 2128 158128 299792
rect 173168 2128 173488 299792
rect 188528 2128 188848 299792
rect 203888 2128 204208 299792
rect 219248 2128 219568 299792
rect 234608 2128 234928 299792
<< obsm4 >>
rect 96843 134675 111648 200293
rect 112128 134675 127008 200293
rect 127488 134675 142368 200293
rect 142848 134675 155789 200293
<< labels >>
rlabel metal2 s 120998 301200 121054 302000 6 adapter_parity
port 1 nsew signal output
rlabel metal2 s 155406 0 155462 800 6 ap_en
port 2 nsew signal output
rlabel metal2 s 17222 0 17278 800 6 clk
port 3 nsew signal input
rlabel metal2 s 51722 0 51778 800 6 clk_en
port 4 nsew signal output
rlabel metal3 s 241200 37680 242000 37800 6 cs_en
port 5 nsew signal output
rlabel metal2 s 24214 301200 24270 302000 6 loopthrough_sel
port 6 nsew signal input
rlabel metal2 s 169390 301200 169446 302000 6 lt_sel_en
port 7 nsew signal output
rlabel metal2 s 72606 301200 72662 302000 6 minion_parity
port 8 nsew signal output
rlabel metal3 s 241200 113160 242000 113280 6 miso_en
port 9 nsew signal output
rlabel metal3 s 241200 188640 242000 188760 6 mosi_en
port 10 nsew signal output
rlabel metal3 s 0 75488 800 75608 6 mp_en
port 11 nsew signal output
rlabel metal2 s 86314 0 86370 800 6 reset
port 12 nsew signal input
rlabel metal2 s 120906 0 120962 800 6 reset_en
port 13 nsew signal output
rlabel metal3 s 241200 264120 242000 264240 6 sclk_en
port 14 nsew signal output
rlabel metal2 s 217782 301200 217838 302000 6 spi_min__cs
port 15 nsew signal input
rlabel metal2 s 189998 0 190054 800 6 spi_min__miso
port 16 nsew signal output
rlabel metal3 s 0 226448 800 226568 6 spi_min__mosi
port 17 nsew signal input
rlabel metal2 s 224590 0 224646 800 6 spi_min__sclk
port 18 nsew signal input
rlabel metal4 s 4208 2128 4528 299792 6 vccd1
port 19 nsew power input
rlabel metal4 s 34928 2128 35248 299792 6 vccd1
port 19 nsew power input
rlabel metal4 s 65648 2128 65968 299792 6 vccd1
port 19 nsew power input
rlabel metal4 s 96368 2128 96688 299792 6 vccd1
port 19 nsew power input
rlabel metal4 s 127088 2128 127408 299792 6 vccd1
port 19 nsew power input
rlabel metal4 s 157808 2128 158128 299792 6 vccd1
port 19 nsew power input
rlabel metal4 s 188528 2128 188848 299792 6 vccd1
port 19 nsew power input
rlabel metal4 s 219248 2128 219568 299792 6 vccd1
port 19 nsew power input
rlabel metal4 s 19568 2128 19888 299792 6 vssd1
port 20 nsew ground input
rlabel metal4 s 50288 2128 50608 299792 6 vssd1
port 20 nsew ground input
rlabel metal4 s 81008 2128 81328 299792 6 vssd1
port 20 nsew ground input
rlabel metal4 s 111728 2128 112048 299792 6 vssd1
port 20 nsew ground input
rlabel metal4 s 142448 2128 142768 299792 6 vssd1
port 20 nsew ground input
rlabel metal4 s 173168 2128 173488 299792 6 vssd1
port 20 nsew ground input
rlabel metal4 s 203888 2128 204208 299792 6 vssd1
port 20 nsew ground input
rlabel metal4 s 234608 2128 234928 299792 6 vssd1
port 20 nsew ground input
<< properties >>
string FIXED_BBOX 0 0 242000 302000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 27191330
string GDS_FILE /home/acm289/ece5745-tapeout/openlane/project-group99/runs/project-group99/results/finishing/grp_99_SPI_TapeOutBlockRTL_32bits_5entries.magic.gds
string GDS_START 512240
<< end >>


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO grp_99_SPI_TapeOutBlockRTL_32bits_5entries
  CLASS BLOCK ;
  FOREIGN grp_99_SPI_TapeOutBlockRTL_32bits_5entries ;
  ORIGIN 0.000 0.000 ;
  SIZE 900.000 BY 900.000 ;
  PIN adapter_parity
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 374.720 900.000 375.320 ;
    END
  END adapter_parity
  PIN ap_en
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 809.690 0.000 809.970 4.000 ;
    END
  END ap_en
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 449.510 0.000 449.790 4.000 ;
    END
  END clk
  PIN clk_en
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 629.830 0.000 630.110 4.000 ;
    END
  END clk_en
  PIN cs_en
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 578.310 896.000 578.590 900.000 ;
    END
  END cs_en
  PIN loopthrough_sel
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 74.840 900.000 75.440 ;
    END
  END loopthrough_sel
  PIN lt_sel_en
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 706.650 896.000 706.930 900.000 ;
    END
  END lt_sel_en
  PIN minion_parity
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 224.440 900.000 225.040 ;
    END
  END minion_parity
  PIN miso_en
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 525.000 900.000 525.600 ;
    END
  END miso_en
  PIN mosi_en
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 835.450 896.000 835.730 900.000 ;
    END
  END mosi_en
  PIN mp_en
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 674.600 900.000 675.200 ;
    END
  END mp_en
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.790 0.000 90.070 4.000 ;
    END
  END reset
  PIN reset_en
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 269.650 0.000 269.930 4.000 ;
    END
  END reset_en
  PIN sclk_en
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 824.880 900.000 825.480 ;
    END
  END sclk_en
  PIN spi_min_cs
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 449.510 896.000 449.790 900.000 ;
    END
  END spi_min_cs
  PIN spi_min_miso
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 192.370 896.000 192.650 900.000 ;
    END
  END spi_min_miso
  PIN spi_min_mosi
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.030 896.000 64.310 900.000 ;
    END
  END spi_min_mosi
  PIN spi_min_sclk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 321.170 896.000 321.450 900.000 ;
    END
  END spi_min_sclk
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 886.960 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 886.960 ;
    END
  END vssd1
  OBS
      LAYER nwell ;
        RECT 5.330 882.585 894.430 885.415 ;
        RECT 5.330 877.145 894.430 879.975 ;
        RECT 5.330 871.705 894.430 874.535 ;
        RECT 5.330 866.265 894.430 869.095 ;
        RECT 5.330 860.825 894.430 863.655 ;
        RECT 5.330 855.385 894.430 858.215 ;
        RECT 5.330 849.945 894.430 852.775 ;
        RECT 5.330 844.505 894.430 847.335 ;
        RECT 5.330 839.065 894.430 841.895 ;
        RECT 5.330 833.625 894.430 836.455 ;
        RECT 5.330 828.185 894.430 831.015 ;
        RECT 5.330 822.745 894.430 825.575 ;
        RECT 5.330 817.305 894.430 820.135 ;
        RECT 5.330 811.865 894.430 814.695 ;
        RECT 5.330 806.425 894.430 809.255 ;
        RECT 5.330 800.985 894.430 803.815 ;
        RECT 5.330 795.545 894.430 798.375 ;
        RECT 5.330 790.105 894.430 792.935 ;
        RECT 5.330 784.665 894.430 787.495 ;
        RECT 5.330 779.225 894.430 782.055 ;
        RECT 5.330 773.785 894.430 776.615 ;
        RECT 5.330 768.345 894.430 771.175 ;
        RECT 5.330 762.905 894.430 765.735 ;
        RECT 5.330 757.465 894.430 760.295 ;
        RECT 5.330 752.025 894.430 754.855 ;
        RECT 5.330 746.585 894.430 749.415 ;
        RECT 5.330 741.145 894.430 743.975 ;
        RECT 5.330 735.705 894.430 738.535 ;
        RECT 5.330 730.265 894.430 733.095 ;
        RECT 5.330 724.825 894.430 727.655 ;
        RECT 5.330 719.385 894.430 722.215 ;
        RECT 5.330 713.945 894.430 716.775 ;
        RECT 5.330 708.505 894.430 711.335 ;
        RECT 5.330 703.065 894.430 705.895 ;
        RECT 5.330 697.625 894.430 700.455 ;
        RECT 5.330 692.185 894.430 695.015 ;
        RECT 5.330 686.745 894.430 689.575 ;
        RECT 5.330 681.305 894.430 684.135 ;
        RECT 5.330 675.865 894.430 678.695 ;
        RECT 5.330 670.425 894.430 673.255 ;
        RECT 5.330 664.985 894.430 667.815 ;
        RECT 5.330 659.545 894.430 662.375 ;
        RECT 5.330 654.105 894.430 656.935 ;
        RECT 5.330 648.665 894.430 651.495 ;
        RECT 5.330 643.225 894.430 646.055 ;
        RECT 5.330 637.785 894.430 640.615 ;
        RECT 5.330 632.345 894.430 635.175 ;
        RECT 5.330 626.905 894.430 629.735 ;
        RECT 5.330 621.465 894.430 624.295 ;
        RECT 5.330 616.025 894.430 618.855 ;
        RECT 5.330 610.585 894.430 613.415 ;
        RECT 5.330 605.145 894.430 607.975 ;
        RECT 5.330 599.705 894.430 602.535 ;
        RECT 5.330 594.265 894.430 597.095 ;
        RECT 5.330 588.825 894.430 591.655 ;
        RECT 5.330 583.385 894.430 586.215 ;
        RECT 5.330 577.945 894.430 580.775 ;
        RECT 5.330 572.505 894.430 575.335 ;
        RECT 5.330 567.065 894.430 569.895 ;
        RECT 5.330 561.625 894.430 564.455 ;
        RECT 5.330 556.185 894.430 559.015 ;
        RECT 5.330 550.745 894.430 553.575 ;
        RECT 5.330 545.305 894.430 548.135 ;
        RECT 5.330 539.865 894.430 542.695 ;
        RECT 5.330 534.425 894.430 537.255 ;
        RECT 5.330 528.985 894.430 531.815 ;
        RECT 5.330 523.545 894.430 526.375 ;
        RECT 5.330 518.105 894.430 520.935 ;
        RECT 5.330 512.665 894.430 515.495 ;
        RECT 5.330 507.225 894.430 510.055 ;
        RECT 5.330 501.785 894.430 504.615 ;
        RECT 5.330 496.345 894.430 499.175 ;
        RECT 5.330 490.905 894.430 493.735 ;
        RECT 5.330 485.465 894.430 488.295 ;
        RECT 5.330 480.025 894.430 482.855 ;
        RECT 5.330 474.585 894.430 477.415 ;
        RECT 5.330 469.145 894.430 471.975 ;
        RECT 5.330 463.705 894.430 466.535 ;
        RECT 5.330 458.265 894.430 461.095 ;
        RECT 5.330 452.825 894.430 455.655 ;
        RECT 5.330 447.385 894.430 450.215 ;
        RECT 5.330 441.945 894.430 444.775 ;
        RECT 5.330 436.505 894.430 439.335 ;
        RECT 5.330 431.065 894.430 433.895 ;
        RECT 5.330 425.625 894.430 428.455 ;
        RECT 5.330 420.185 894.430 423.015 ;
        RECT 5.330 414.745 894.430 417.575 ;
        RECT 5.330 409.305 894.430 412.135 ;
        RECT 5.330 403.865 894.430 406.695 ;
        RECT 5.330 398.425 894.430 401.255 ;
        RECT 5.330 392.985 894.430 395.815 ;
        RECT 5.330 387.545 894.430 390.375 ;
        RECT 5.330 382.105 894.430 384.935 ;
        RECT 5.330 376.665 894.430 379.495 ;
        RECT 5.330 371.225 894.430 374.055 ;
        RECT 5.330 365.785 894.430 368.615 ;
        RECT 5.330 360.345 894.430 363.175 ;
        RECT 5.330 354.905 894.430 357.735 ;
        RECT 5.330 349.465 894.430 352.295 ;
        RECT 5.330 344.025 894.430 346.855 ;
        RECT 5.330 338.585 894.430 341.415 ;
        RECT 5.330 333.145 894.430 335.975 ;
        RECT 5.330 327.705 894.430 330.535 ;
        RECT 5.330 322.265 894.430 325.095 ;
        RECT 5.330 316.825 894.430 319.655 ;
        RECT 5.330 311.385 894.430 314.215 ;
        RECT 5.330 305.945 894.430 308.775 ;
        RECT 5.330 300.505 894.430 303.335 ;
        RECT 5.330 295.065 894.430 297.895 ;
        RECT 5.330 289.625 894.430 292.455 ;
        RECT 5.330 284.185 894.430 287.015 ;
        RECT 5.330 278.745 894.430 281.575 ;
        RECT 5.330 273.305 894.430 276.135 ;
        RECT 5.330 267.865 894.430 270.695 ;
        RECT 5.330 262.425 894.430 265.255 ;
        RECT 5.330 256.985 894.430 259.815 ;
        RECT 5.330 251.545 894.430 254.375 ;
        RECT 5.330 246.105 894.430 248.935 ;
        RECT 5.330 240.665 894.430 243.495 ;
        RECT 5.330 235.225 894.430 238.055 ;
        RECT 5.330 229.785 894.430 232.615 ;
        RECT 5.330 224.345 894.430 227.175 ;
        RECT 5.330 218.905 894.430 221.735 ;
        RECT 5.330 213.465 894.430 216.295 ;
        RECT 5.330 208.025 894.430 210.855 ;
        RECT 5.330 202.585 894.430 205.415 ;
        RECT 5.330 197.145 894.430 199.975 ;
        RECT 5.330 191.705 894.430 194.535 ;
        RECT 5.330 186.265 894.430 189.095 ;
        RECT 5.330 180.825 894.430 183.655 ;
        RECT 5.330 175.385 894.430 178.215 ;
        RECT 5.330 169.945 894.430 172.775 ;
        RECT 5.330 164.505 894.430 167.335 ;
        RECT 5.330 159.065 894.430 161.895 ;
        RECT 5.330 153.625 894.430 156.455 ;
        RECT 5.330 148.185 894.430 151.015 ;
        RECT 5.330 142.745 894.430 145.575 ;
        RECT 5.330 137.305 894.430 140.135 ;
        RECT 5.330 131.865 894.430 134.695 ;
        RECT 5.330 126.425 894.430 129.255 ;
        RECT 5.330 120.985 894.430 123.815 ;
        RECT 5.330 115.545 894.430 118.375 ;
        RECT 5.330 110.105 894.430 112.935 ;
        RECT 5.330 104.665 894.430 107.495 ;
        RECT 5.330 99.225 894.430 102.055 ;
        RECT 5.330 93.785 894.430 96.615 ;
        RECT 5.330 88.345 894.430 91.175 ;
        RECT 5.330 82.905 894.430 85.735 ;
        RECT 5.330 77.465 894.430 80.295 ;
        RECT 5.330 72.025 894.430 74.855 ;
        RECT 5.330 66.585 894.430 69.415 ;
        RECT 5.330 61.145 894.430 63.975 ;
        RECT 5.330 55.705 894.430 58.535 ;
        RECT 5.330 50.265 894.430 53.095 ;
        RECT 5.330 44.825 894.430 47.655 ;
        RECT 5.330 39.385 894.430 42.215 ;
        RECT 5.330 33.945 894.430 36.775 ;
        RECT 5.330 28.505 894.430 31.335 ;
        RECT 5.330 23.065 894.430 25.895 ;
        RECT 5.330 17.625 894.430 20.455 ;
        RECT 5.330 12.185 894.430 15.015 ;
      LAYER li1 ;
        RECT 5.520 10.795 894.240 886.805 ;
      LAYER met1 ;
        RECT 5.520 10.640 894.240 886.960 ;
      LAYER met2 ;
        RECT 21.070 895.720 63.750 896.650 ;
        RECT 64.590 895.720 192.090 896.650 ;
        RECT 192.930 895.720 320.890 896.650 ;
        RECT 321.730 895.720 449.230 896.650 ;
        RECT 450.070 895.720 578.030 896.650 ;
        RECT 578.870 895.720 706.370 896.650 ;
        RECT 707.210 895.720 835.170 896.650 ;
        RECT 836.010 895.720 890.930 896.650 ;
        RECT 21.070 4.280 890.930 895.720 ;
        RECT 21.070 4.000 89.510 4.280 ;
        RECT 90.350 4.000 269.370 4.280 ;
        RECT 270.210 4.000 449.230 4.280 ;
        RECT 450.070 4.000 629.550 4.280 ;
        RECT 630.390 4.000 809.410 4.280 ;
        RECT 810.250 4.000 890.930 4.280 ;
      LAYER met3 ;
        RECT 21.040 825.880 896.000 886.885 ;
        RECT 21.040 824.480 895.600 825.880 ;
        RECT 21.040 675.600 896.000 824.480 ;
        RECT 21.040 674.200 895.600 675.600 ;
        RECT 21.040 526.000 896.000 674.200 ;
        RECT 21.040 524.600 895.600 526.000 ;
        RECT 21.040 375.720 896.000 524.600 ;
        RECT 21.040 374.320 895.600 375.720 ;
        RECT 21.040 225.440 896.000 374.320 ;
        RECT 21.040 224.040 895.600 225.440 ;
        RECT 21.040 75.840 896.000 224.040 ;
        RECT 21.040 74.440 895.600 75.840 ;
        RECT 21.040 10.715 896.000 74.440 ;
      LAYER met4 ;
        RECT 548.615 16.495 558.240 579.865 ;
        RECT 560.640 16.495 602.305 579.865 ;
  END
END grp_99_SPI_TapeOutBlockRTL_32bits_5entries
END LIBRARY


magic
tech sky130A
magscale 1 2
timestamp 1655438056
<< obsli1 >>
rect 1104 2159 138828 137649
<< obsm1 >>
rect 1104 2128 138828 137680
<< metal2 >>
rect 14002 139200 14058 140000
rect 41970 139200 42026 140000
rect 69938 139200 69994 140000
rect 97998 139200 98054 140000
rect 125966 139200 126022 140000
rect 17498 0 17554 800
rect 52458 0 52514 800
rect 87510 0 87566 800
rect 122470 0 122526 800
<< obsm2 >>
rect 1398 139144 13946 139346
rect 14114 139144 41914 139346
rect 42082 139144 69882 139346
rect 70050 139144 97942 139346
rect 98110 139144 125910 139346
rect 126078 139144 138166 139346
rect 1398 856 138166 139144
rect 1398 800 17442 856
rect 17610 800 52402 856
rect 52570 800 87454 856
rect 87622 800 122414 856
rect 122582 800 138166 856
<< metal3 >>
rect 0 128120 800 128240
rect 139200 116560 140000 116680
rect 0 104864 800 104984
rect 0 81472 800 81592
rect 139200 69912 140000 70032
rect 0 58216 800 58336
rect 0 34824 800 34944
rect 139200 23264 140000 23384
rect 0 11568 800 11688
<< obsm3 >>
rect 800 128320 139200 137665
rect 880 128040 139200 128320
rect 800 116760 139200 128040
rect 800 116480 139120 116760
rect 800 105064 139200 116480
rect 880 104784 139200 105064
rect 800 81672 139200 104784
rect 880 81392 139200 81672
rect 800 70112 139200 81392
rect 800 69832 139120 70112
rect 800 58416 139200 69832
rect 880 58136 139200 58416
rect 800 35024 139200 58136
rect 880 34744 139200 35024
rect 800 23464 139200 34744
rect 800 23184 139120 23464
rect 800 11768 139200 23184
rect 880 11488 139200 11768
rect 800 2143 139200 11488
<< metal4 >>
rect 4208 2128 4528 137680
rect 19568 2128 19888 137680
rect 34928 2128 35248 137680
rect 50288 2128 50608 137680
rect 65648 2128 65968 137680
rect 81008 2128 81328 137680
rect 96368 2128 96688 137680
rect 111728 2128 112048 137680
rect 127088 2128 127408 137680
<< obsm4 >>
rect 11651 23563 19488 135285
rect 19968 23563 34848 135285
rect 35328 23563 50208 135285
rect 50688 23563 65568 135285
rect 66048 23563 80928 135285
rect 81408 23563 96288 135285
rect 96768 23563 111648 135285
rect 112128 23563 127008 135285
rect 127488 23563 137941 135285
<< labels >>
rlabel metal2 s 87510 0 87566 800 6 adapter_parity
port 1 nsew signal output
rlabel metal2 s 125966 139200 126022 140000 6 ap_en
port 2 nsew signal output
rlabel metal2 s 14002 139200 14058 140000 6 clk
port 3 nsew signal input
rlabel metal2 s 41970 139200 42026 140000 6 clk_en
port 4 nsew signal output
rlabel metal2 s 122470 0 122526 800 6 cs_en
port 5 nsew signal output
rlabel metal3 s 0 58216 800 58336 6 loopthrough_sel
port 6 nsew signal input
rlabel metal3 s 0 104864 800 104984 6 lt_sel_en
port 7 nsew signal output
rlabel metal3 s 0 81472 800 81592 6 minion_parity
port 8 nsew signal output
rlabel metal3 s 139200 23264 140000 23384 6 miso_en
port 9 nsew signal output
rlabel metal3 s 0 128120 800 128240 6 mosi_en
port 10 nsew signal output
rlabel metal3 s 139200 69912 140000 70032 6 mp_en
port 11 nsew signal output
rlabel metal2 s 69938 139200 69994 140000 6 reset
port 12 nsew signal input
rlabel metal2 s 97998 139200 98054 140000 6 reset_en
port 13 nsew signal output
rlabel metal3 s 139200 116560 140000 116680 6 sclk_en
port 14 nsew signal output
rlabel metal2 s 52458 0 52514 800 6 spi_min_cs
port 15 nsew signal input
rlabel metal3 s 0 11568 800 11688 6 spi_min_miso
port 16 nsew signal output
rlabel metal3 s 0 34824 800 34944 6 spi_min_mosi
port 17 nsew signal input
rlabel metal2 s 17498 0 17554 800 6 spi_min_sclk
port 18 nsew signal input
rlabel metal4 s 4208 2128 4528 137680 6 vccd1
port 19 nsew power input
rlabel metal4 s 34928 2128 35248 137680 6 vccd1
port 19 nsew power input
rlabel metal4 s 65648 2128 65968 137680 6 vccd1
port 19 nsew power input
rlabel metal4 s 96368 2128 96688 137680 6 vccd1
port 19 nsew power input
rlabel metal4 s 127088 2128 127408 137680 6 vccd1
port 19 nsew power input
rlabel metal4 s 19568 2128 19888 137680 6 vssd1
port 20 nsew ground input
rlabel metal4 s 50288 2128 50608 137680 6 vssd1
port 20 nsew ground input
rlabel metal4 s 81008 2128 81328 137680 6 vssd1
port 20 nsew ground input
rlabel metal4 s 111728 2128 112048 137680 6 vssd1
port 20 nsew ground input
<< properties >>
string FIXED_BBOX 0 0 140000 140000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 31617820
string GDS_FILE /home/acm289/ece5745-tapeout/openlane/project-group17/runs/project-group17/results/finishing/grp_17_SPI_TapeOutBlockRTL_32bits_5entries.magic.gds
string GDS_START 1410736
<< end >>


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO grp_15_SPI_TapeOutBlockRTL_32bits_5entries
  CLASS BLOCK ;
  FOREIGN grp_15_SPI_TapeOutBlockRTL_32bits_5entries ;
  ORIGIN 0.000 0.000 ;
  SIZE 900.000 BY 900.000 ;
  PIN adapter_parity
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 74.840 900.000 75.440 ;
    END
  END adapter_parity
  PIN ap_en
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 693.640 900.000 694.240 ;
    END
  END ap_en
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 508.850 896.000 509.130 900.000 ;
    END
  END clk
  PIN clk_en
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 582.910 0.000 583.190 4.000 ;
    END
  END clk_en
  PIN cs_en
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 822.840 4.000 823.440 ;
    END
  END cs_en
  PIN loopthrough_sel
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 315.650 896.000 315.930 900.000 ;
    END
  END loopthrough_sel
  PIN lt_sel_en
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END lt_sel_en
  PIN minion_parity
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 898.470 896.000 898.750 900.000 ;
    END
  END minion_parity
  PIN miso_en
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 779.330 0.000 779.610 4.000 ;
    END
  END miso_en
  PIN mosi_en
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.290 0.000 193.570 4.000 ;
    END
  END mosi_en
  PIN mp_en
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 204.040 4.000 204.640 ;
    END
  END mp_en
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 486.240 900.000 486.840 ;
    END
  END reset
  PIN reset_en
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 411.440 4.000 412.040 ;
    END
  END reset_en
  PIN sclk_en
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 705.270 896.000 705.550 900.000 ;
    END
  END sclk_en
  PIN spi_min_cs
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 389.710 0.000 389.990 4.000 ;
    END
  END spi_min_cs
  PIN spi_min_miso
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 615.440 4.000 616.040 ;
    END
  END spi_min_miso
  PIN spi_min_mosi
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.230 896.000 119.510 900.000 ;
    END
  END spi_min_mosi
  PIN spi_min_sclk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 282.240 900.000 282.840 ;
    END
  END spi_min_sclk
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 886.960 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 886.960 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 894.240 886.805 ;
      LAYER met1 ;
        RECT 0.070 10.640 898.770 886.960 ;
      LAYER met2 ;
        RECT 0.100 895.720 118.950 896.650 ;
        RECT 119.790 895.720 315.370 896.650 ;
        RECT 316.210 895.720 508.570 896.650 ;
        RECT 509.410 895.720 704.990 896.650 ;
        RECT 705.830 895.720 898.190 896.650 ;
        RECT 0.100 4.280 898.740 895.720 ;
        RECT 0.650 4.000 193.010 4.280 ;
        RECT 193.850 4.000 389.430 4.280 ;
        RECT 390.270 4.000 582.630 4.280 ;
        RECT 583.470 4.000 779.050 4.280 ;
        RECT 779.890 4.000 898.740 4.280 ;
      LAYER met3 ;
        RECT 4.000 823.840 896.000 886.885 ;
        RECT 4.400 822.440 896.000 823.840 ;
        RECT 4.000 694.640 896.000 822.440 ;
        RECT 4.000 693.240 895.600 694.640 ;
        RECT 4.000 616.440 896.000 693.240 ;
        RECT 4.400 615.040 896.000 616.440 ;
        RECT 4.000 487.240 896.000 615.040 ;
        RECT 4.000 485.840 895.600 487.240 ;
        RECT 4.000 412.440 896.000 485.840 ;
        RECT 4.400 411.040 896.000 412.440 ;
        RECT 4.000 283.240 896.000 411.040 ;
        RECT 4.000 281.840 895.600 283.240 ;
        RECT 4.000 205.040 896.000 281.840 ;
        RECT 4.400 203.640 896.000 205.040 ;
        RECT 4.000 75.840 896.000 203.640 ;
        RECT 4.000 74.440 895.600 75.840 ;
        RECT 4.000 10.715 896.000 74.440 ;
      LAYER met4 ;
        RECT 326.895 329.975 327.840 659.425 ;
        RECT 330.240 329.975 404.640 659.425 ;
        RECT 407.040 329.975 481.440 659.425 ;
        RECT 483.840 329.975 558.240 659.425 ;
        RECT 560.640 329.975 635.040 659.425 ;
        RECT 637.440 329.975 684.185 659.425 ;
  END
END grp_15_SPI_TapeOutBlockRTL_32bits_5entries
END LIBRARY


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO grp_99_SPI_TapeOutBlockRTL_32bits_5entries
  CLASS BLOCK ;
  FOREIGN grp_99_SPI_TapeOutBlockRTL_32bits_5entries ;
  ORIGIN 0.000 0.000 ;
  SIZE 700.000 BY 700.000 ;
  PIN adapter_parity
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 582.800 700.000 583.400 ;
    END
  END adapter_parity
  PIN ap_en
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 116.320 4.000 116.920 ;
    END
  END ap_en
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 291.270 0.000 291.550 4.000 ;
    END
  END clk
  PIN clk_en
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 408.110 0.000 408.390 4.000 ;
    END
  END clk_en
  PIN cs_en
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 349.560 4.000 350.160 ;
    END
  END cs_en
  PIN loopthrough_sel
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 116.320 700.000 116.920 ;
    END
  END loopthrough_sel
  PIN lt_sel_en
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 524.490 696.000 524.770 700.000 ;
    END
  END lt_sel_en
  PIN minion_parity
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 349.560 700.000 350.160 ;
    END
  END minion_parity
  PIN miso_en
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 582.800 4.000 583.400 ;
    END
  END miso_en
  PIN mosi_en
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 524.490 0.000 524.770 4.000 ;
    END
  END mosi_en
  PIN mp_en
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 641.330 696.000 641.610 700.000 ;
    END
  END mp_en
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.050 0.000 58.330 4.000 ;
    END
  END reset
  PIN reset_en
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 174.430 0.000 174.710 4.000 ;
    END
  END reset_en
  PIN sclk_en
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 641.330 0.000 641.610 4.000 ;
    END
  END sclk_en
  PIN spi_min_cs
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 408.110 696.000 408.390 700.000 ;
    END
  END spi_min_cs
  PIN spi_min_miso
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 174.430 696.000 174.710 700.000 ;
    END
  END spi_min_miso
  PIN spi_min_mosi
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.050 696.000 58.330 700.000 ;
    END
  END spi_min_mosi
  PIN spi_min_sclk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 291.270 696.000 291.550 700.000 ;
    END
  END spi_min_sclk
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 688.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 688.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 688.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 688.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 688.400 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 688.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 688.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 688.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 688.400 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 694.140 688.245 ;
      LAYER met1 ;
        RECT 5.520 10.640 694.140 688.400 ;
      LAYER met2 ;
        RECT 6.990 695.720 57.770 696.730 ;
        RECT 58.610 695.720 174.150 696.730 ;
        RECT 174.990 695.720 290.990 696.730 ;
        RECT 291.830 695.720 407.830 696.730 ;
        RECT 408.670 695.720 524.210 696.730 ;
        RECT 525.050 695.720 641.050 696.730 ;
        RECT 641.890 695.720 690.830 696.730 ;
        RECT 6.990 4.280 690.830 695.720 ;
        RECT 6.990 4.000 57.770 4.280 ;
        RECT 58.610 4.000 174.150 4.280 ;
        RECT 174.990 4.000 290.990 4.280 ;
        RECT 291.830 4.000 407.830 4.280 ;
        RECT 408.670 4.000 524.210 4.280 ;
        RECT 525.050 4.000 641.050 4.280 ;
        RECT 641.890 4.000 690.830 4.280 ;
      LAYER met3 ;
        RECT 4.000 583.800 696.000 688.325 ;
        RECT 4.400 582.400 695.600 583.800 ;
        RECT 4.000 350.560 696.000 582.400 ;
        RECT 4.400 349.160 695.600 350.560 ;
        RECT 4.000 117.320 696.000 349.160 ;
        RECT 4.400 115.920 695.600 117.320 ;
        RECT 4.000 10.715 696.000 115.920 ;
      LAYER met4 ;
        RECT 389.455 118.495 404.640 586.665 ;
        RECT 407.040 118.495 454.185 586.665 ;
  END
END grp_99_SPI_TapeOutBlockRTL_32bits_5entries
END LIBRARY


magic
tech sky130A
magscale 1 2
timestamp 1654199528
<< nwell >>
rect 1066 299461 240894 299782
rect 1066 298373 240894 298939
rect 1066 297285 240894 297851
rect 1066 296197 240894 296763
rect 1066 295109 240894 295675
rect 1066 294021 240894 294587
rect 1066 292933 240894 293499
rect 1066 291845 240894 292411
rect 1066 290757 240894 291323
rect 1066 289669 240894 290235
rect 1066 288581 240894 289147
rect 1066 287493 240894 288059
rect 1066 286405 240894 286971
rect 1066 285317 240894 285883
rect 1066 284229 240894 284795
rect 1066 283141 240894 283707
rect 1066 282053 240894 282619
rect 1066 280965 240894 281531
rect 1066 279877 240894 280443
rect 1066 278789 240894 279355
rect 1066 277701 240894 278267
rect 1066 276613 240894 277179
rect 1066 275525 240894 276091
rect 1066 274437 240894 275003
rect 1066 273349 240894 273915
rect 1066 272261 240894 272827
rect 1066 271173 240894 271739
rect 1066 270085 240894 270651
rect 1066 268997 240894 269563
rect 1066 267909 240894 268475
rect 1066 266821 240894 267387
rect 1066 265733 240894 266299
rect 1066 264645 240894 265211
rect 1066 263557 240894 264123
rect 1066 262469 240894 263035
rect 1066 261381 240894 261947
rect 1066 260293 240894 260859
rect 1066 259205 240894 259771
rect 1066 258117 240894 258683
rect 1066 257029 240894 257595
rect 1066 255941 240894 256507
rect 1066 254853 240894 255419
rect 1066 253765 240894 254331
rect 1066 252677 240894 253243
rect 1066 251589 240894 252155
rect 1066 250501 240894 251067
rect 1066 249413 240894 249979
rect 1066 248325 240894 248891
rect 1066 247237 240894 247803
rect 1066 246149 240894 246715
rect 1066 245061 240894 245627
rect 1066 243973 240894 244539
rect 1066 242885 240894 243451
rect 1066 241797 240894 242363
rect 1066 240709 240894 241275
rect 1066 239621 240894 240187
rect 1066 238533 240894 239099
rect 1066 237445 240894 238011
rect 1066 236357 240894 236923
rect 1066 235269 240894 235835
rect 1066 234181 240894 234747
rect 1066 233093 240894 233659
rect 1066 232005 240894 232571
rect 1066 230917 240894 231483
rect 1066 229829 240894 230395
rect 1066 228741 240894 229307
rect 1066 227653 240894 228219
rect 1066 226565 240894 227131
rect 1066 225477 240894 226043
rect 1066 224389 240894 224955
rect 1066 223301 240894 223867
rect 1066 222213 240894 222779
rect 1066 221125 240894 221691
rect 1066 220037 240894 220603
rect 1066 218949 240894 219515
rect 1066 217861 240894 218427
rect 1066 216773 240894 217339
rect 1066 215685 240894 216251
rect 1066 214597 240894 215163
rect 1066 213509 240894 214075
rect 1066 212421 240894 212987
rect 1066 211333 240894 211899
rect 1066 210245 240894 210811
rect 1066 209157 240894 209723
rect 1066 208069 240894 208635
rect 1066 206981 240894 207547
rect 1066 205893 240894 206459
rect 1066 204805 240894 205371
rect 1066 203717 240894 204283
rect 1066 202629 240894 203195
rect 1066 201541 240894 202107
rect 1066 200453 240894 201019
rect 1066 199365 240894 199931
rect 1066 198277 240894 198843
rect 1066 197189 240894 197755
rect 1066 196101 240894 196667
rect 1066 195013 240894 195579
rect 1066 193925 240894 194491
rect 1066 192837 240894 193403
rect 1066 191749 240894 192315
rect 1066 190661 240894 191227
rect 1066 189573 240894 190139
rect 1066 188485 240894 189051
rect 1066 187397 240894 187963
rect 1066 186309 240894 186875
rect 1066 185221 240894 185787
rect 1066 184133 240894 184699
rect 1066 183045 240894 183611
rect 1066 181957 240894 182523
rect 1066 180869 240894 181435
rect 1066 179781 240894 180347
rect 1066 178693 240894 179259
rect 1066 177605 240894 178171
rect 1066 176517 240894 177083
rect 1066 175429 240894 175995
rect 1066 174341 240894 174907
rect 1066 173253 240894 173819
rect 1066 172165 240894 172731
rect 1066 171077 240894 171643
rect 1066 169989 240894 170555
rect 1066 168901 240894 169467
rect 1066 167813 240894 168379
rect 1066 166725 240894 167291
rect 1066 165637 240894 166203
rect 1066 164549 240894 165115
rect 1066 163461 240894 164027
rect 1066 162373 240894 162939
rect 1066 161285 240894 161851
rect 1066 160197 240894 160763
rect 1066 159109 240894 159675
rect 1066 158021 240894 158587
rect 1066 156933 240894 157499
rect 1066 155845 240894 156411
rect 1066 154757 240894 155323
rect 1066 153669 240894 154235
rect 1066 152581 240894 153147
rect 1066 151493 240894 152059
rect 1066 150405 240894 150971
rect 1066 149317 240894 149883
rect 1066 148229 240894 148795
rect 1066 147141 240894 147707
rect 1066 146053 240894 146619
rect 1066 144965 240894 145531
rect 1066 143877 240894 144443
rect 1066 142789 240894 143355
rect 1066 141701 240894 142267
rect 1066 140613 240894 141179
rect 1066 139525 240894 140091
rect 1066 138437 240894 139003
rect 1066 137349 240894 137915
rect 1066 136261 240894 136827
rect 1066 135173 240894 135739
rect 1066 134085 240894 134651
rect 1066 132997 240894 133563
rect 1066 131909 240894 132475
rect 1066 130821 240894 131387
rect 1066 129733 240894 130299
rect 1066 128645 240894 129211
rect 1066 127557 240894 128123
rect 1066 126469 240894 127035
rect 1066 125381 240894 125947
rect 1066 124293 240894 124859
rect 1066 123205 240894 123771
rect 1066 122117 240894 122683
rect 1066 121029 240894 121595
rect 1066 119941 240894 120507
rect 1066 118853 240894 119419
rect 1066 117765 240894 118331
rect 1066 116677 240894 117243
rect 1066 115589 240894 116155
rect 1066 114501 240894 115067
rect 1066 113413 240894 113979
rect 1066 112325 240894 112891
rect 1066 111237 240894 111803
rect 1066 110149 240894 110715
rect 1066 109061 240894 109627
rect 1066 107973 240894 108539
rect 1066 106885 240894 107451
rect 1066 105797 240894 106363
rect 1066 104709 240894 105275
rect 1066 103621 240894 104187
rect 1066 102533 240894 103099
rect 1066 101445 240894 102011
rect 1066 100357 240894 100923
rect 1066 99269 240894 99835
rect 1066 98181 240894 98747
rect 1066 97093 240894 97659
rect 1066 96005 240894 96571
rect 1066 94917 240894 95483
rect 1066 93829 240894 94395
rect 1066 92741 240894 93307
rect 1066 91653 240894 92219
rect 1066 90565 240894 91131
rect 1066 89477 240894 90043
rect 1066 88389 240894 88955
rect 1066 87301 240894 87867
rect 1066 86213 240894 86779
rect 1066 85125 240894 85691
rect 1066 84037 240894 84603
rect 1066 82949 240894 83515
rect 1066 81861 240894 82427
rect 1066 80773 240894 81339
rect 1066 79685 240894 80251
rect 1066 78597 240894 79163
rect 1066 77509 240894 78075
rect 1066 76421 240894 76987
rect 1066 75333 240894 75899
rect 1066 74245 240894 74811
rect 1066 73157 240894 73723
rect 1066 72069 240894 72635
rect 1066 70981 240894 71547
rect 1066 69893 240894 70459
rect 1066 68805 240894 69371
rect 1066 67717 240894 68283
rect 1066 66629 240894 67195
rect 1066 65541 240894 66107
rect 1066 64453 240894 65019
rect 1066 63365 240894 63931
rect 1066 62277 240894 62843
rect 1066 61189 240894 61755
rect 1066 60101 240894 60667
rect 1066 59013 240894 59579
rect 1066 57925 240894 58491
rect 1066 56837 240894 57403
rect 1066 55749 240894 56315
rect 1066 54661 240894 55227
rect 1066 53573 240894 54139
rect 1066 52485 240894 53051
rect 1066 51397 240894 51963
rect 1066 50309 240894 50875
rect 1066 49221 240894 49787
rect 1066 48133 240894 48699
rect 1066 47045 240894 47611
rect 1066 45957 240894 46523
rect 1066 44869 240894 45435
rect 1066 43781 240894 44347
rect 1066 42693 240894 43259
rect 1066 41605 240894 42171
rect 1066 40517 240894 41083
rect 1066 39429 240894 39995
rect 1066 38341 240894 38907
rect 1066 37253 240894 37819
rect 1066 36165 240894 36731
rect 1066 35077 240894 35643
rect 1066 33989 240894 34555
rect 1066 32901 240894 33467
rect 1066 31813 240894 32379
rect 1066 30725 240894 31291
rect 1066 29637 240894 30203
rect 1066 28549 240894 29115
rect 1066 27461 240894 28027
rect 1066 26373 240894 26939
rect 1066 25285 240894 25851
rect 1066 24197 240894 24763
rect 1066 23109 240894 23675
rect 1066 22021 240894 22587
rect 1066 20933 240894 21499
rect 1066 19845 240894 20411
rect 1066 18757 240894 19323
rect 1066 17669 240894 18235
rect 1066 16581 240894 17147
rect 1066 15493 240894 16059
rect 1066 14405 240894 14971
rect 1066 13317 240894 13883
rect 1066 12229 240894 12795
rect 1066 11141 240894 11707
rect 1066 10053 240894 10619
rect 1066 8965 240894 9531
rect 1066 7877 240894 8443
rect 1066 6789 240894 7355
rect 1066 5701 240894 6267
rect 1066 4613 240894 5179
rect 1066 3525 240894 4091
rect 1066 2437 240894 3003
<< obsli1 >>
rect 1104 2159 240856 299761
<< obsm1 >>
rect 1104 2128 240856 299792
<< metal2 >>
rect 30194 301200 30250 302000
rect 90638 301200 90694 302000
rect 151174 301200 151230 302000
rect 211618 301200 211674 302000
rect 30194 0 30250 800
rect 90638 0 90694 800
rect 151174 0 151230 800
rect 211618 0 211674 800
<< obsm2 >>
rect 4214 301144 30138 301322
rect 30306 301144 90582 301322
rect 90750 301144 151118 301322
rect 151286 301144 211562 301322
rect 211730 301144 240194 301322
rect 4214 856 240194 301144
rect 4214 734 30138 856
rect 30306 734 90582 856
rect 90750 734 151118 856
rect 151286 734 211562 856
rect 211730 734 240194 856
<< metal3 >>
rect 241200 150968 242000 151088
<< obsm3 >>
rect 4208 151168 241200 299777
rect 4208 150888 241120 151168
rect 4208 2143 241200 150888
<< metal4 >>
rect 4208 2128 4528 299792
rect 19568 2128 19888 299792
rect 34928 2128 35248 299792
rect 50288 2128 50608 299792
rect 65648 2128 65968 299792
rect 81008 2128 81328 299792
rect 96368 2128 96688 299792
rect 111728 2128 112048 299792
rect 127088 2128 127408 299792
rect 142448 2128 142768 299792
rect 157808 2128 158128 299792
rect 173168 2128 173488 299792
rect 188528 2128 188848 299792
rect 203888 2128 204208 299792
rect 219248 2128 219568 299792
rect 234608 2128 234928 299792
<< obsm4 >>
rect 127571 107475 142368 190501
rect 142848 107475 157728 190501
rect 158208 107475 173088 190501
rect 173568 107475 186149 190501
<< labels >>
rlabel metal2 s 151174 301200 151230 302000 6 adapter_parity
port 1 nsew signal output
rlabel metal2 s 30194 0 30250 800 6 clk
port 2 nsew signal input
rlabel metal2 s 30194 301200 30250 302000 6 loopthrough_sel
port 3 nsew signal input
rlabel metal2 s 90638 301200 90694 302000 6 minion_parity
port 4 nsew signal output
rlabel metal2 s 90638 0 90694 800 6 reset
port 5 nsew signal input
rlabel metal2 s 151174 0 151230 800 6 spi_min__cs
port 6 nsew signal input
rlabel metal2 s 211618 0 211674 800 6 spi_min__miso
port 7 nsew signal output
rlabel metal2 s 211618 301200 211674 302000 6 spi_min__mosi
port 8 nsew signal input
rlabel metal3 s 241200 150968 242000 151088 6 spi_min__sclk
port 9 nsew signal input
rlabel metal4 s 4208 2128 4528 299792 6 vccd1
port 10 nsew power input
rlabel metal4 s 34928 2128 35248 299792 6 vccd1
port 10 nsew power input
rlabel metal4 s 65648 2128 65968 299792 6 vccd1
port 10 nsew power input
rlabel metal4 s 96368 2128 96688 299792 6 vccd1
port 10 nsew power input
rlabel metal4 s 127088 2128 127408 299792 6 vccd1
port 10 nsew power input
rlabel metal4 s 157808 2128 158128 299792 6 vccd1
port 10 nsew power input
rlabel metal4 s 188528 2128 188848 299792 6 vccd1
port 10 nsew power input
rlabel metal4 s 219248 2128 219568 299792 6 vccd1
port 10 nsew power input
rlabel metal4 s 19568 2128 19888 299792 6 vssd1
port 11 nsew ground input
rlabel metal4 s 50288 2128 50608 299792 6 vssd1
port 11 nsew ground input
rlabel metal4 s 81008 2128 81328 299792 6 vssd1
port 11 nsew ground input
rlabel metal4 s 111728 2128 112048 299792 6 vssd1
port 11 nsew ground input
rlabel metal4 s 142448 2128 142768 299792 6 vssd1
port 11 nsew ground input
rlabel metal4 s 173168 2128 173488 299792 6 vssd1
port 11 nsew ground input
rlabel metal4 s 203888 2128 204208 299792 6 vssd1
port 11 nsew ground input
rlabel metal4 s 234608 2128 234928 299792 6 vssd1
port 11 nsew ground input
<< properties >>
string FIXED_BBOX 0 0 242000 302000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 27345858
string GDS_FILE /home/acm289/ece5745-tapeout/openlane/project-group99/runs/project-group99/results/finishing/grp_99_SPI_TapeOutBlockRTL_32bits_5entries.magic.gds
string GDS_START 486174
<< end >>


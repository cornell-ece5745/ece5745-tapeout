magic
tech sky130A
magscale 1 2
timestamp 1655402207
<< obsli1 >>
rect 1104 2159 240856 299761
<< obsm1 >>
rect 1104 2128 240856 299792
<< metal2 >>
rect 30194 301200 30250 302000
rect 90638 301200 90694 302000
rect 151174 301200 151230 302000
rect 211618 301200 211674 302000
rect 24214 0 24270 800
rect 72606 0 72662 800
rect 120998 0 121054 800
rect 169390 0 169446 800
rect 217782 0 217838 800
<< obsm2 >>
rect 1398 301144 30138 301322
rect 30306 301144 90582 301322
rect 90750 301144 151118 301322
rect 151286 301144 211562 301322
rect 211730 301144 240194 301322
rect 1398 856 240194 301144
rect 1398 734 24158 856
rect 24326 734 72550 856
rect 72718 734 120942 856
rect 121110 734 169334 856
rect 169502 734 217726 856
rect 217894 734 240194 856
<< metal3 >>
rect 241200 276768 242000 276888
rect 0 251608 800 251728
rect 241200 226448 242000 226568
rect 241200 176128 242000 176248
rect 0 150968 800 151088
rect 241200 125808 242000 125928
rect 241200 75488 242000 75608
rect 0 50328 800 50448
rect 241200 25168 242000 25288
<< obsm3 >>
rect 800 276968 241200 299777
rect 800 276688 241120 276968
rect 800 251808 241200 276688
rect 880 251528 241200 251808
rect 800 226648 241200 251528
rect 800 226368 241120 226648
rect 800 176328 241200 226368
rect 800 176048 241120 176328
rect 800 151168 241200 176048
rect 880 150888 241200 151168
rect 800 126008 241200 150888
rect 800 125728 241120 126008
rect 800 75688 241200 125728
rect 800 75408 241120 75688
rect 800 50528 241200 75408
rect 880 50248 241200 50528
rect 800 25368 241200 50248
rect 800 25088 241120 25368
rect 800 2143 241200 25088
<< metal4 >>
rect 4208 2128 4528 299792
rect 19568 2128 19888 299792
rect 34928 2128 35248 299792
rect 50288 2128 50608 299792
rect 65648 2128 65968 299792
rect 81008 2128 81328 299792
rect 96368 2128 96688 299792
rect 111728 2128 112048 299792
rect 127088 2128 127408 299792
rect 142448 2128 142768 299792
rect 157808 2128 158128 299792
rect 173168 2128 173488 299792
rect 188528 2128 188848 299792
rect 203888 2128 204208 299792
rect 219248 2128 219568 299792
rect 234608 2128 234928 299792
<< obsm4 >>
rect 118555 147731 127008 225997
rect 127488 147731 142368 225997
rect 142848 147731 157728 225997
rect 158208 147731 173088 225997
rect 173568 147731 188357 225997
<< labels >>
rlabel metal2 s 151174 301200 151230 302000 6 adapter_parity
port 1 nsew signal output
rlabel metal3 s 0 50328 800 50448 6 ap_en
port 2 nsew signal output
rlabel metal2 s 24214 0 24270 800 6 clk
port 3 nsew signal input
rlabel metal2 s 72606 0 72662 800 6 clk_en
port 4 nsew signal output
rlabel metal3 s 0 150968 800 151088 6 cs_en
port 5 nsew signal output
rlabel metal2 s 30194 301200 30250 302000 6 loopthrough_sel
port 6 nsew signal input
rlabel metal3 s 241200 226448 242000 226568 6 lt_sel_en
port 7 nsew signal output
rlabel metal2 s 90638 301200 90694 302000 6 minion_parity
port 8 nsew signal output
rlabel metal2 s 217782 0 217838 800 6 miso_en
port 9 nsew signal output
rlabel metal3 s 0 251608 800 251728 6 mosi_en
port 10 nsew signal output
rlabel metal2 s 211618 301200 211674 302000 6 mp_en
port 11 nsew signal output
rlabel metal2 s 120998 0 121054 800 6 reset
port 12 nsew signal input
rlabel metal2 s 169390 0 169446 800 6 reset_en
port 13 nsew signal output
rlabel metal3 s 241200 276768 242000 276888 6 sclk_en
port 14 nsew signal output
rlabel metal3 s 241200 25168 242000 25288 6 spi_min_cs
port 15 nsew signal input
rlabel metal3 s 241200 75488 242000 75608 6 spi_min_miso
port 16 nsew signal output
rlabel metal3 s 241200 125808 242000 125928 6 spi_min_mosi
port 17 nsew signal input
rlabel metal3 s 241200 176128 242000 176248 6 spi_min_sclk
port 18 nsew signal input
rlabel metal4 s 4208 2128 4528 299792 6 vccd1
port 19 nsew power input
rlabel metal4 s 34928 2128 35248 299792 6 vccd1
port 19 nsew power input
rlabel metal4 s 65648 2128 65968 299792 6 vccd1
port 19 nsew power input
rlabel metal4 s 96368 2128 96688 299792 6 vccd1
port 19 nsew power input
rlabel metal4 s 127088 2128 127408 299792 6 vccd1
port 19 nsew power input
rlabel metal4 s 157808 2128 158128 299792 6 vccd1
port 19 nsew power input
rlabel metal4 s 188528 2128 188848 299792 6 vccd1
port 19 nsew power input
rlabel metal4 s 219248 2128 219568 299792 6 vccd1
port 19 nsew power input
rlabel metal4 s 19568 2128 19888 299792 6 vssd1
port 20 nsew ground input
rlabel metal4 s 50288 2128 50608 299792 6 vssd1
port 20 nsew ground input
rlabel metal4 s 81008 2128 81328 299792 6 vssd1
port 20 nsew ground input
rlabel metal4 s 111728 2128 112048 299792 6 vssd1
port 20 nsew ground input
rlabel metal4 s 142448 2128 142768 299792 6 vssd1
port 20 nsew ground input
rlabel metal4 s 173168 2128 173488 299792 6 vssd1
port 20 nsew ground input
rlabel metal4 s 203888 2128 204208 299792 6 vssd1
port 20 nsew ground input
rlabel metal4 s 234608 2128 234928 299792 6 vssd1
port 20 nsew ground input
<< properties >>
string FIXED_BBOX 0 0 242000 302000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 29340846
string GDS_FILE /home/acm289/ece5745-tapeout/openlane/project-group99/runs/project-group99/results/finishing/grp_99_SPI_TapeOutBlockRTL_32bits_5entries.magic.gds
string GDS_START 625848
<< end >>


magic
tech sky130A
magscale 1 2
timestamp 1655481690
<< nwell >>
rect 1066 176517 178886 177083
rect 1066 175429 178886 175995
rect 1066 174341 178886 174907
rect 1066 173253 178886 173819
rect 1066 172165 178886 172731
rect 1066 171077 178886 171643
rect 1066 169989 178886 170555
rect 1066 168901 178886 169467
rect 1066 167813 178886 168379
rect 1066 166725 178886 167291
rect 1066 165637 178886 166203
rect 1066 164549 178886 165115
rect 1066 163461 178886 164027
rect 1066 162373 178886 162939
rect 1066 161285 178886 161851
rect 1066 160197 178886 160763
rect 1066 159109 178886 159675
rect 1066 158021 178886 158587
rect 1066 156933 178886 157499
rect 1066 155845 178886 156411
rect 1066 154757 178886 155323
rect 1066 153669 178886 154235
rect 1066 152581 178886 153147
rect 1066 151493 178886 152059
rect 1066 150405 178886 150971
rect 1066 149317 178886 149883
rect 1066 148229 178886 148795
rect 1066 147141 178886 147707
rect 1066 146053 178886 146619
rect 1066 144965 178886 145531
rect 1066 143877 178886 144443
rect 1066 142789 178886 143355
rect 1066 141701 178886 142267
rect 1066 140613 178886 141179
rect 1066 139525 178886 140091
rect 1066 138437 178886 139003
rect 1066 137349 178886 137915
rect 1066 136261 178886 136827
rect 1066 135173 178886 135739
rect 1066 134085 178886 134651
rect 1066 132997 178886 133563
rect 1066 131909 178886 132475
rect 1066 130821 178886 131387
rect 1066 129733 178886 130299
rect 1066 128645 178886 129211
rect 1066 127557 178886 128123
rect 1066 126469 178886 127035
rect 1066 125381 178886 125947
rect 1066 124293 178886 124859
rect 1066 123205 178886 123771
rect 1066 122117 178886 122683
rect 1066 121029 178886 121595
rect 1066 119941 178886 120507
rect 1066 118853 178886 119419
rect 1066 117765 178886 118331
rect 1066 116677 178886 117243
rect 1066 115589 178886 116155
rect 1066 114501 178886 115067
rect 1066 113413 178886 113979
rect 1066 112325 178886 112891
rect 1066 111237 178886 111803
rect 1066 110149 178886 110715
rect 1066 109061 178886 109627
rect 1066 107973 178886 108539
rect 1066 106885 178886 107451
rect 1066 105797 178886 106363
rect 1066 104709 178886 105275
rect 1066 103621 178886 104187
rect 1066 102533 178886 103099
rect 1066 101445 178886 102011
rect 1066 100357 178886 100923
rect 1066 99269 178886 99835
rect 1066 98181 178886 98747
rect 1066 97093 178886 97659
rect 1066 96005 178886 96571
rect 1066 94917 178886 95483
rect 1066 93829 178886 94395
rect 1066 92741 178886 93307
rect 1066 91653 178886 92219
rect 1066 90565 178886 91131
rect 1066 89477 178886 90043
rect 1066 88389 178886 88955
rect 1066 87301 178886 87867
rect 1066 86213 178886 86779
rect 1066 85125 178886 85691
rect 1066 84037 178886 84603
rect 1066 82949 178886 83515
rect 1066 81861 178886 82427
rect 1066 80773 178886 81339
rect 1066 79685 178886 80251
rect 1066 78597 178886 79163
rect 1066 77509 178886 78075
rect 1066 76421 178886 76987
rect 1066 75333 178886 75899
rect 1066 74245 178886 74811
rect 1066 73157 178886 73723
rect 1066 72069 178886 72635
rect 1066 70981 178886 71547
rect 1066 69893 178886 70459
rect 1066 68805 178886 69371
rect 1066 67717 178886 68283
rect 1066 66629 178886 67195
rect 1066 65541 178886 66107
rect 1066 64453 178886 65019
rect 1066 63365 178886 63931
rect 1066 62277 178886 62843
rect 1066 61189 178886 61755
rect 1066 60101 178886 60667
rect 1066 59013 178886 59579
rect 1066 57925 178886 58491
rect 1066 56837 178886 57403
rect 1066 55749 178886 56315
rect 1066 54661 178886 55227
rect 1066 53573 178886 54139
rect 1066 52485 178886 53051
rect 1066 51397 178886 51963
rect 1066 50309 178886 50875
rect 1066 49221 178886 49787
rect 1066 48133 178886 48699
rect 1066 47045 178886 47611
rect 1066 45957 178886 46523
rect 1066 44869 178886 45435
rect 1066 43781 178886 44347
rect 1066 42693 178886 43259
rect 1066 41605 178886 42171
rect 1066 40517 178886 41083
rect 1066 39429 178886 39995
rect 1066 38341 178886 38907
rect 1066 37253 178886 37819
rect 1066 36165 178886 36731
rect 1066 35077 178886 35643
rect 1066 33989 178886 34555
rect 1066 32901 178886 33467
rect 1066 31813 178886 32379
rect 1066 30725 178886 31291
rect 1066 29637 178886 30203
rect 1066 28549 178886 29115
rect 1066 27461 178886 28027
rect 1066 26373 178886 26939
rect 1066 25285 178886 25851
rect 1066 24197 178886 24763
rect 1066 23109 178886 23675
rect 1066 22021 178886 22587
rect 1066 20933 178886 21499
rect 1066 19845 178886 20411
rect 1066 18757 178886 19323
rect 1066 17669 178886 18235
rect 1066 16581 178886 17147
rect 1066 15493 178886 16059
rect 1066 14405 178886 14971
rect 1066 13317 178886 13883
rect 1066 12229 178886 12795
rect 1066 11141 178886 11707
rect 1066 10053 178886 10619
rect 1066 8965 178886 9531
rect 1066 7877 178886 8443
rect 1066 6789 178886 7355
rect 1066 5701 178886 6267
rect 1066 4613 178886 5179
rect 1066 3525 178886 4091
rect 1066 2437 178886 3003
<< obsli1 >>
rect 1104 2159 178848 177361
<< obsm1 >>
rect 1104 2128 178848 177392
<< metal2 >>
rect 12806 179200 12862 180000
rect 38474 179200 38530 180000
rect 64234 179200 64290 180000
rect 89902 179200 89958 180000
rect 115662 179200 115718 180000
rect 141330 179200 141386 180000
rect 167090 179200 167146 180000
rect 17958 0 18014 800
rect 53930 0 53986 800
rect 89902 0 89958 800
rect 125966 0 126022 800
rect 161938 0 161994 800
<< obsm2 >>
rect 4214 179144 12750 179330
rect 12918 179144 38418 179330
rect 38586 179144 64178 179330
rect 64346 179144 89846 179330
rect 90014 179144 115606 179330
rect 115774 179144 141274 179330
rect 141442 179144 167034 179330
rect 167202 179144 178186 179330
rect 4214 856 178186 179144
rect 4214 800 17902 856
rect 18070 800 53874 856
rect 54042 800 89846 856
rect 90014 800 125910 856
rect 126078 800 161882 856
rect 162050 800 178186 856
<< metal3 >>
rect 179200 164976 180000 165096
rect 179200 134920 180000 135040
rect 179200 105000 180000 105120
rect 179200 74944 180000 75064
rect 179200 44888 180000 45008
rect 179200 14968 180000 15088
<< obsm3 >>
rect 4208 165176 179200 177377
rect 4208 164896 179120 165176
rect 4208 135120 179200 164896
rect 4208 134840 179120 135120
rect 4208 105200 179200 134840
rect 4208 104920 179120 105200
rect 4208 75144 179200 104920
rect 4208 74864 179120 75144
rect 4208 45088 179200 74864
rect 4208 44808 179120 45088
rect 4208 15168 179200 44808
rect 4208 14888 179120 15168
rect 4208 2143 179200 14888
<< metal4 >>
rect 4208 2128 4528 177392
rect 19568 2128 19888 177392
rect 34928 2128 35248 177392
rect 50288 2128 50608 177392
rect 65648 2128 65968 177392
rect 81008 2128 81328 177392
rect 96368 2128 96688 177392
rect 111728 2128 112048 177392
rect 127088 2128 127408 177392
rect 142448 2128 142768 177392
rect 157808 2128 158128 177392
rect 173168 2128 173488 177392
<< obsm4 >>
rect 109723 3299 111648 115973
rect 112128 3299 120461 115973
<< labels >>
rlabel metal3 s 179200 74944 180000 75064 6 adapter_parity
port 1 nsew signal output
rlabel metal2 s 161938 0 161994 800 6 ap_en
port 2 nsew signal output
rlabel metal2 s 89902 0 89958 800 6 clk
port 3 nsew signal input
rlabel metal2 s 125966 0 126022 800 6 clk_en
port 4 nsew signal output
rlabel metal2 s 115662 179200 115718 180000 6 cs_en
port 5 nsew signal output
rlabel metal3 s 179200 14968 180000 15088 6 loopthrough_sel
port 6 nsew signal input
rlabel metal2 s 141330 179200 141386 180000 6 lt_sel_en
port 7 nsew signal output
rlabel metal3 s 179200 44888 180000 45008 6 minion_parity
port 8 nsew signal output
rlabel metal3 s 179200 105000 180000 105120 6 miso_en
port 9 nsew signal output
rlabel metal2 s 167090 179200 167146 180000 6 mosi_en
port 10 nsew signal output
rlabel metal3 s 179200 134920 180000 135040 6 mp_en
port 11 nsew signal output
rlabel metal2 s 17958 0 18014 800 6 reset
port 12 nsew signal input
rlabel metal2 s 53930 0 53986 800 6 reset_en
port 13 nsew signal output
rlabel metal3 s 179200 164976 180000 165096 6 sclk_en
port 14 nsew signal output
rlabel metal2 s 89902 179200 89958 180000 6 spi_min_cs
port 15 nsew signal input
rlabel metal2 s 38474 179200 38530 180000 6 spi_min_miso
port 16 nsew signal output
rlabel metal2 s 12806 179200 12862 180000 6 spi_min_mosi
port 17 nsew signal input
rlabel metal2 s 64234 179200 64290 180000 6 spi_min_sclk
port 18 nsew signal input
rlabel metal4 s 4208 2128 4528 177392 6 vccd1
port 19 nsew power input
rlabel metal4 s 34928 2128 35248 177392 6 vccd1
port 19 nsew power input
rlabel metal4 s 65648 2128 65968 177392 6 vccd1
port 19 nsew power input
rlabel metal4 s 96368 2128 96688 177392 6 vccd1
port 19 nsew power input
rlabel metal4 s 127088 2128 127408 177392 6 vccd1
port 19 nsew power input
rlabel metal4 s 157808 2128 158128 177392 6 vccd1
port 19 nsew power input
rlabel metal4 s 19568 2128 19888 177392 6 vssd1
port 20 nsew ground input
rlabel metal4 s 50288 2128 50608 177392 6 vssd1
port 20 nsew ground input
rlabel metal4 s 81008 2128 81328 177392 6 vssd1
port 20 nsew ground input
rlabel metal4 s 111728 2128 112048 177392 6 vssd1
port 20 nsew ground input
rlabel metal4 s 142448 2128 142768 177392 6 vssd1
port 20 nsew ground input
rlabel metal4 s 173168 2128 173488 177392 6 vssd1
port 20 nsew ground input
<< properties >>
string FIXED_BBOX 0 0 180000 180000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 15252614
string GDS_FILE /home/acm289/ece5745-tapeout/openlane/project-group99/runs/project-group99/results/finishing/grp_99_SPI_TapeOutBlockRTL_32bits_5entries.magic.gds
string GDS_START 666340
<< end >>


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO grp_99_SPI_TapeOutBlockRTL_32bits_5entries
  CLASS BLOCK ;
  FOREIGN grp_99_SPI_TapeOutBlockRTL_32bits_5entries ;
  ORIGIN 0.000 0.000 ;
  SIZE 1210.000 BY 1510.000 ;
  PIN adapter_parity
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1007.950 1506.000 1008.230 1510.000 ;
    END
  END adapter_parity
  PIN ap_en
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1206.000 970.400 1210.000 971.000 ;
    END
  END ap_en
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.110 0.000 86.390 4.000 ;
    END
  END clk
  PIN clk_en
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 258.610 0.000 258.890 4.000 ;
    END
  END clk_en
  PIN cs_en
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1206.000 107.480 1210.000 108.080 ;
    END
  END cs_en
  PIN loopthrough_sel
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 201.570 1506.000 201.850 1510.000 ;
    END
  END loopthrough_sel
  PIN lt_sel_en
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 754.840 4.000 755.440 ;
    END
  END lt_sel_en
  PIN minion_parity
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 604.530 1506.000 604.810 1510.000 ;
    END
  END minion_parity
  PIN miso_en
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1206.000 323.040 1210.000 323.640 ;
    END
  END miso_en
  PIN mosi_en
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1206.000 538.600 1210.000 539.200 ;
    END
  END mosi_en
  PIN mp_en
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1206.000 1185.960 1210.000 1186.560 ;
    END
  END mp_en
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 431.570 0.000 431.850 4.000 ;
    END
  END reset
  PIN reset_en
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 604.530 0.000 604.810 4.000 ;
    END
  END reset_en
  PIN sclk_en
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1206.000 754.160 1210.000 754.760 ;
    END
  END sclk_en
  PIN spi_min__cs
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 777.030 0.000 777.310 4.000 ;
    END
  END spi_min__cs
  PIN spi_min__miso
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1206.000 1401.520 1210.000 1402.120 ;
    END
  END spi_min__miso
  PIN spi_min__mosi
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 949.990 0.000 950.270 4.000 ;
    END
  END spi_min__mosi
  PIN spi_min__sclk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1122.950 0.000 1123.230 4.000 ;
    END
  END spi_min__sclk
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 1498.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 1498.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 1498.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 1498.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 1498.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 1498.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 942.640 10.640 944.240 1498.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 1096.240 10.640 1097.840 1498.960 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 1498.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 1498.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 1498.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 1498.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 1498.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 1498.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 1019.440 10.640 1021.040 1498.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 1173.040 10.640 1174.640 1498.960 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 1204.280 1498.805 ;
      LAYER met1 ;
        RECT 5.520 10.640 1204.280 1498.960 ;
      LAYER met2 ;
        RECT 6.990 1505.720 201.290 1506.610 ;
        RECT 202.130 1505.720 604.250 1506.610 ;
        RECT 605.090 1505.720 1007.670 1506.610 ;
        RECT 1008.510 1505.720 1200.970 1506.610 ;
        RECT 6.990 4.280 1200.970 1505.720 ;
        RECT 6.990 3.670 85.830 4.280 ;
        RECT 86.670 3.670 258.330 4.280 ;
        RECT 259.170 3.670 431.290 4.280 ;
        RECT 432.130 3.670 604.250 4.280 ;
        RECT 605.090 3.670 776.750 4.280 ;
        RECT 777.590 3.670 949.710 4.280 ;
        RECT 950.550 3.670 1122.670 4.280 ;
        RECT 1123.510 3.670 1200.970 4.280 ;
      LAYER met3 ;
        RECT 4.000 1402.520 1206.000 1498.885 ;
        RECT 4.000 1401.120 1205.600 1402.520 ;
        RECT 4.000 1186.960 1206.000 1401.120 ;
        RECT 4.000 1185.560 1205.600 1186.960 ;
        RECT 4.000 971.400 1206.000 1185.560 ;
        RECT 4.000 970.000 1205.600 971.400 ;
        RECT 4.000 755.840 1206.000 970.000 ;
        RECT 4.400 755.160 1206.000 755.840 ;
        RECT 4.400 754.440 1205.600 755.160 ;
        RECT 4.000 753.760 1205.600 754.440 ;
        RECT 4.000 539.600 1206.000 753.760 ;
        RECT 4.000 538.200 1205.600 539.600 ;
        RECT 4.000 324.040 1206.000 538.200 ;
        RECT 4.000 322.640 1205.600 324.040 ;
        RECT 4.000 108.480 1206.000 322.640 ;
        RECT 4.000 107.080 1205.600 108.480 ;
        RECT 4.000 10.715 1206.000 107.080 ;
      LAYER met4 ;
        RECT 668.215 631.895 711.840 945.705 ;
        RECT 714.240 631.895 788.640 945.705 ;
        RECT 791.040 631.895 865.440 945.705 ;
        RECT 867.840 631.895 942.240 945.705 ;
        RECT 944.640 631.895 1019.040 945.705 ;
        RECT 1021.440 631.895 1046.665 945.705 ;
  END
END grp_99_SPI_TapeOutBlockRTL_32bits_5entries
END LIBRARY


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO grp_99_SPI_TapeOutBlockRTL_32bits_5entries
  CLASS BLOCK ;
  FOREIGN grp_99_SPI_TapeOutBlockRTL_32bits_5entries ;
  ORIGIN 0.000 0.000 ;
  SIZE 1210.000 BY 1510.000 ;
  PIN adapter_parity
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 755.870 1506.000 756.150 1510.000 ;
    END
  END adapter_parity
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.970 0.000 151.250 4.000 ;
    END
  END clk
  PIN loopthrough_sel
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.970 1506.000 151.250 1510.000 ;
    END
  END loopthrough_sel
  PIN minion_parity
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 453.190 1506.000 453.470 1510.000 ;
    END
  END minion_parity
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 453.190 0.000 453.470 4.000 ;
    END
  END reset
  PIN spi_min__cs
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 755.870 0.000 756.150 4.000 ;
    END
  END spi_min__cs
  PIN spi_min__miso
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1058.090 0.000 1058.370 4.000 ;
    END
  END spi_min__miso
  PIN spi_min__mosi
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1058.090 1506.000 1058.370 1510.000 ;
    END
  END spi_min__mosi
  PIN spi_min__sclk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1206.000 754.840 1210.000 755.440 ;
    END
  END spi_min__sclk
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 1498.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 1498.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 1498.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 1498.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 1498.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 1498.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 942.640 10.640 944.240 1498.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 1096.240 10.640 1097.840 1498.960 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 1498.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 1498.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 1498.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 1498.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 1498.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 1498.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 1019.440 10.640 1021.040 1498.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 1173.040 10.640 1174.640 1498.960 ;
    END
  END vssd1
  OBS
      LAYER nwell ;
        RECT 5.330 1497.305 1204.470 1498.910 ;
        RECT 5.330 1491.865 1204.470 1494.695 ;
        RECT 5.330 1486.425 1204.470 1489.255 ;
        RECT 5.330 1480.985 1204.470 1483.815 ;
        RECT 5.330 1475.545 1204.470 1478.375 ;
        RECT 5.330 1470.105 1204.470 1472.935 ;
        RECT 5.330 1464.665 1204.470 1467.495 ;
        RECT 5.330 1459.225 1204.470 1462.055 ;
        RECT 5.330 1453.785 1204.470 1456.615 ;
        RECT 5.330 1448.345 1204.470 1451.175 ;
        RECT 5.330 1442.905 1204.470 1445.735 ;
        RECT 5.330 1437.465 1204.470 1440.295 ;
        RECT 5.330 1432.025 1204.470 1434.855 ;
        RECT 5.330 1426.585 1204.470 1429.415 ;
        RECT 5.330 1421.145 1204.470 1423.975 ;
        RECT 5.330 1415.705 1204.470 1418.535 ;
        RECT 5.330 1410.265 1204.470 1413.095 ;
        RECT 5.330 1404.825 1204.470 1407.655 ;
        RECT 5.330 1399.385 1204.470 1402.215 ;
        RECT 5.330 1393.945 1204.470 1396.775 ;
        RECT 5.330 1388.505 1204.470 1391.335 ;
        RECT 5.330 1383.065 1204.470 1385.895 ;
        RECT 5.330 1377.625 1204.470 1380.455 ;
        RECT 5.330 1372.185 1204.470 1375.015 ;
        RECT 5.330 1366.745 1204.470 1369.575 ;
        RECT 5.330 1361.305 1204.470 1364.135 ;
        RECT 5.330 1355.865 1204.470 1358.695 ;
        RECT 5.330 1350.425 1204.470 1353.255 ;
        RECT 5.330 1344.985 1204.470 1347.815 ;
        RECT 5.330 1339.545 1204.470 1342.375 ;
        RECT 5.330 1334.105 1204.470 1336.935 ;
        RECT 5.330 1328.665 1204.470 1331.495 ;
        RECT 5.330 1323.225 1204.470 1326.055 ;
        RECT 5.330 1317.785 1204.470 1320.615 ;
        RECT 5.330 1312.345 1204.470 1315.175 ;
        RECT 5.330 1306.905 1204.470 1309.735 ;
        RECT 5.330 1301.465 1204.470 1304.295 ;
        RECT 5.330 1296.025 1204.470 1298.855 ;
        RECT 5.330 1290.585 1204.470 1293.415 ;
        RECT 5.330 1285.145 1204.470 1287.975 ;
        RECT 5.330 1279.705 1204.470 1282.535 ;
        RECT 5.330 1274.265 1204.470 1277.095 ;
        RECT 5.330 1268.825 1204.470 1271.655 ;
        RECT 5.330 1263.385 1204.470 1266.215 ;
        RECT 5.330 1257.945 1204.470 1260.775 ;
        RECT 5.330 1252.505 1204.470 1255.335 ;
        RECT 5.330 1247.065 1204.470 1249.895 ;
        RECT 5.330 1241.625 1204.470 1244.455 ;
        RECT 5.330 1236.185 1204.470 1239.015 ;
        RECT 5.330 1230.745 1204.470 1233.575 ;
        RECT 5.330 1225.305 1204.470 1228.135 ;
        RECT 5.330 1219.865 1204.470 1222.695 ;
        RECT 5.330 1214.425 1204.470 1217.255 ;
        RECT 5.330 1208.985 1204.470 1211.815 ;
        RECT 5.330 1203.545 1204.470 1206.375 ;
        RECT 5.330 1198.105 1204.470 1200.935 ;
        RECT 5.330 1192.665 1204.470 1195.495 ;
        RECT 5.330 1187.225 1204.470 1190.055 ;
        RECT 5.330 1181.785 1204.470 1184.615 ;
        RECT 5.330 1176.345 1204.470 1179.175 ;
        RECT 5.330 1170.905 1204.470 1173.735 ;
        RECT 5.330 1165.465 1204.470 1168.295 ;
        RECT 5.330 1160.025 1204.470 1162.855 ;
        RECT 5.330 1154.585 1204.470 1157.415 ;
        RECT 5.330 1149.145 1204.470 1151.975 ;
        RECT 5.330 1143.705 1204.470 1146.535 ;
        RECT 5.330 1138.265 1204.470 1141.095 ;
        RECT 5.330 1132.825 1204.470 1135.655 ;
        RECT 5.330 1127.385 1204.470 1130.215 ;
        RECT 5.330 1121.945 1204.470 1124.775 ;
        RECT 5.330 1116.505 1204.470 1119.335 ;
        RECT 5.330 1111.065 1204.470 1113.895 ;
        RECT 5.330 1105.625 1204.470 1108.455 ;
        RECT 5.330 1100.185 1204.470 1103.015 ;
        RECT 5.330 1094.745 1204.470 1097.575 ;
        RECT 5.330 1089.305 1204.470 1092.135 ;
        RECT 5.330 1083.865 1204.470 1086.695 ;
        RECT 5.330 1078.425 1204.470 1081.255 ;
        RECT 5.330 1072.985 1204.470 1075.815 ;
        RECT 5.330 1067.545 1204.470 1070.375 ;
        RECT 5.330 1062.105 1204.470 1064.935 ;
        RECT 5.330 1056.665 1204.470 1059.495 ;
        RECT 5.330 1051.225 1204.470 1054.055 ;
        RECT 5.330 1045.785 1204.470 1048.615 ;
        RECT 5.330 1040.345 1204.470 1043.175 ;
        RECT 5.330 1034.905 1204.470 1037.735 ;
        RECT 5.330 1029.465 1204.470 1032.295 ;
        RECT 5.330 1024.025 1204.470 1026.855 ;
        RECT 5.330 1018.585 1204.470 1021.415 ;
        RECT 5.330 1013.145 1204.470 1015.975 ;
        RECT 5.330 1007.705 1204.470 1010.535 ;
        RECT 5.330 1002.265 1204.470 1005.095 ;
        RECT 5.330 996.825 1204.470 999.655 ;
        RECT 5.330 991.385 1204.470 994.215 ;
        RECT 5.330 985.945 1204.470 988.775 ;
        RECT 5.330 980.505 1204.470 983.335 ;
        RECT 5.330 975.065 1204.470 977.895 ;
        RECT 5.330 969.625 1204.470 972.455 ;
        RECT 5.330 964.185 1204.470 967.015 ;
        RECT 5.330 958.745 1204.470 961.575 ;
        RECT 5.330 953.305 1204.470 956.135 ;
        RECT 5.330 947.865 1204.470 950.695 ;
        RECT 5.330 942.425 1204.470 945.255 ;
        RECT 5.330 936.985 1204.470 939.815 ;
        RECT 5.330 931.545 1204.470 934.375 ;
        RECT 5.330 926.105 1204.470 928.935 ;
        RECT 5.330 920.665 1204.470 923.495 ;
        RECT 5.330 915.225 1204.470 918.055 ;
        RECT 5.330 909.785 1204.470 912.615 ;
        RECT 5.330 904.345 1204.470 907.175 ;
        RECT 5.330 898.905 1204.470 901.735 ;
        RECT 5.330 893.465 1204.470 896.295 ;
        RECT 5.330 888.025 1204.470 890.855 ;
        RECT 5.330 882.585 1204.470 885.415 ;
        RECT 5.330 877.145 1204.470 879.975 ;
        RECT 5.330 871.705 1204.470 874.535 ;
        RECT 5.330 866.265 1204.470 869.095 ;
        RECT 5.330 860.825 1204.470 863.655 ;
        RECT 5.330 855.385 1204.470 858.215 ;
        RECT 5.330 849.945 1204.470 852.775 ;
        RECT 5.330 844.505 1204.470 847.335 ;
        RECT 5.330 839.065 1204.470 841.895 ;
        RECT 5.330 833.625 1204.470 836.455 ;
        RECT 5.330 828.185 1204.470 831.015 ;
        RECT 5.330 822.745 1204.470 825.575 ;
        RECT 5.330 817.305 1204.470 820.135 ;
        RECT 5.330 811.865 1204.470 814.695 ;
        RECT 5.330 806.425 1204.470 809.255 ;
        RECT 5.330 800.985 1204.470 803.815 ;
        RECT 5.330 795.545 1204.470 798.375 ;
        RECT 5.330 790.105 1204.470 792.935 ;
        RECT 5.330 784.665 1204.470 787.495 ;
        RECT 5.330 779.225 1204.470 782.055 ;
        RECT 5.330 773.785 1204.470 776.615 ;
        RECT 5.330 768.345 1204.470 771.175 ;
        RECT 5.330 762.905 1204.470 765.735 ;
        RECT 5.330 757.465 1204.470 760.295 ;
        RECT 5.330 752.025 1204.470 754.855 ;
        RECT 5.330 746.585 1204.470 749.415 ;
        RECT 5.330 741.145 1204.470 743.975 ;
        RECT 5.330 735.705 1204.470 738.535 ;
        RECT 5.330 730.265 1204.470 733.095 ;
        RECT 5.330 724.825 1204.470 727.655 ;
        RECT 5.330 719.385 1204.470 722.215 ;
        RECT 5.330 713.945 1204.470 716.775 ;
        RECT 5.330 708.505 1204.470 711.335 ;
        RECT 5.330 703.065 1204.470 705.895 ;
        RECT 5.330 697.625 1204.470 700.455 ;
        RECT 5.330 692.185 1204.470 695.015 ;
        RECT 5.330 686.745 1204.470 689.575 ;
        RECT 5.330 681.305 1204.470 684.135 ;
        RECT 5.330 675.865 1204.470 678.695 ;
        RECT 5.330 670.425 1204.470 673.255 ;
        RECT 5.330 664.985 1204.470 667.815 ;
        RECT 5.330 659.545 1204.470 662.375 ;
        RECT 5.330 654.105 1204.470 656.935 ;
        RECT 5.330 648.665 1204.470 651.495 ;
        RECT 5.330 643.225 1204.470 646.055 ;
        RECT 5.330 637.785 1204.470 640.615 ;
        RECT 5.330 632.345 1204.470 635.175 ;
        RECT 5.330 626.905 1204.470 629.735 ;
        RECT 5.330 621.465 1204.470 624.295 ;
        RECT 5.330 616.025 1204.470 618.855 ;
        RECT 5.330 610.585 1204.470 613.415 ;
        RECT 5.330 605.145 1204.470 607.975 ;
        RECT 5.330 599.705 1204.470 602.535 ;
        RECT 5.330 594.265 1204.470 597.095 ;
        RECT 5.330 588.825 1204.470 591.655 ;
        RECT 5.330 583.385 1204.470 586.215 ;
        RECT 5.330 577.945 1204.470 580.775 ;
        RECT 5.330 572.505 1204.470 575.335 ;
        RECT 5.330 567.065 1204.470 569.895 ;
        RECT 5.330 561.625 1204.470 564.455 ;
        RECT 5.330 556.185 1204.470 559.015 ;
        RECT 5.330 550.745 1204.470 553.575 ;
        RECT 5.330 545.305 1204.470 548.135 ;
        RECT 5.330 539.865 1204.470 542.695 ;
        RECT 5.330 534.425 1204.470 537.255 ;
        RECT 5.330 528.985 1204.470 531.815 ;
        RECT 5.330 523.545 1204.470 526.375 ;
        RECT 5.330 518.105 1204.470 520.935 ;
        RECT 5.330 512.665 1204.470 515.495 ;
        RECT 5.330 507.225 1204.470 510.055 ;
        RECT 5.330 501.785 1204.470 504.615 ;
        RECT 5.330 496.345 1204.470 499.175 ;
        RECT 5.330 490.905 1204.470 493.735 ;
        RECT 5.330 485.465 1204.470 488.295 ;
        RECT 5.330 480.025 1204.470 482.855 ;
        RECT 5.330 474.585 1204.470 477.415 ;
        RECT 5.330 469.145 1204.470 471.975 ;
        RECT 5.330 463.705 1204.470 466.535 ;
        RECT 5.330 458.265 1204.470 461.095 ;
        RECT 5.330 452.825 1204.470 455.655 ;
        RECT 5.330 447.385 1204.470 450.215 ;
        RECT 5.330 441.945 1204.470 444.775 ;
        RECT 5.330 436.505 1204.470 439.335 ;
        RECT 5.330 431.065 1204.470 433.895 ;
        RECT 5.330 425.625 1204.470 428.455 ;
        RECT 5.330 420.185 1204.470 423.015 ;
        RECT 5.330 414.745 1204.470 417.575 ;
        RECT 5.330 409.305 1204.470 412.135 ;
        RECT 5.330 403.865 1204.470 406.695 ;
        RECT 5.330 398.425 1204.470 401.255 ;
        RECT 5.330 392.985 1204.470 395.815 ;
        RECT 5.330 387.545 1204.470 390.375 ;
        RECT 5.330 382.105 1204.470 384.935 ;
        RECT 5.330 376.665 1204.470 379.495 ;
        RECT 5.330 371.225 1204.470 374.055 ;
        RECT 5.330 365.785 1204.470 368.615 ;
        RECT 5.330 360.345 1204.470 363.175 ;
        RECT 5.330 354.905 1204.470 357.735 ;
        RECT 5.330 349.465 1204.470 352.295 ;
        RECT 5.330 344.025 1204.470 346.855 ;
        RECT 5.330 338.585 1204.470 341.415 ;
        RECT 5.330 333.145 1204.470 335.975 ;
        RECT 5.330 327.705 1204.470 330.535 ;
        RECT 5.330 322.265 1204.470 325.095 ;
        RECT 5.330 316.825 1204.470 319.655 ;
        RECT 5.330 311.385 1204.470 314.215 ;
        RECT 5.330 305.945 1204.470 308.775 ;
        RECT 5.330 300.505 1204.470 303.335 ;
        RECT 5.330 295.065 1204.470 297.895 ;
        RECT 5.330 289.625 1204.470 292.455 ;
        RECT 5.330 284.185 1204.470 287.015 ;
        RECT 5.330 278.745 1204.470 281.575 ;
        RECT 5.330 273.305 1204.470 276.135 ;
        RECT 5.330 267.865 1204.470 270.695 ;
        RECT 5.330 262.425 1204.470 265.255 ;
        RECT 5.330 256.985 1204.470 259.815 ;
        RECT 5.330 251.545 1204.470 254.375 ;
        RECT 5.330 246.105 1204.470 248.935 ;
        RECT 5.330 240.665 1204.470 243.495 ;
        RECT 5.330 235.225 1204.470 238.055 ;
        RECT 5.330 229.785 1204.470 232.615 ;
        RECT 5.330 224.345 1204.470 227.175 ;
        RECT 5.330 218.905 1204.470 221.735 ;
        RECT 5.330 213.465 1204.470 216.295 ;
        RECT 5.330 208.025 1204.470 210.855 ;
        RECT 5.330 202.585 1204.470 205.415 ;
        RECT 5.330 197.145 1204.470 199.975 ;
        RECT 5.330 191.705 1204.470 194.535 ;
        RECT 5.330 186.265 1204.470 189.095 ;
        RECT 5.330 180.825 1204.470 183.655 ;
        RECT 5.330 175.385 1204.470 178.215 ;
        RECT 5.330 169.945 1204.470 172.775 ;
        RECT 5.330 164.505 1204.470 167.335 ;
        RECT 5.330 159.065 1204.470 161.895 ;
        RECT 5.330 153.625 1204.470 156.455 ;
        RECT 5.330 148.185 1204.470 151.015 ;
        RECT 5.330 142.745 1204.470 145.575 ;
        RECT 5.330 137.305 1204.470 140.135 ;
        RECT 5.330 131.865 1204.470 134.695 ;
        RECT 5.330 126.425 1204.470 129.255 ;
        RECT 5.330 120.985 1204.470 123.815 ;
        RECT 5.330 115.545 1204.470 118.375 ;
        RECT 5.330 110.105 1204.470 112.935 ;
        RECT 5.330 104.665 1204.470 107.495 ;
        RECT 5.330 99.225 1204.470 102.055 ;
        RECT 5.330 93.785 1204.470 96.615 ;
        RECT 5.330 88.345 1204.470 91.175 ;
        RECT 5.330 82.905 1204.470 85.735 ;
        RECT 5.330 77.465 1204.470 80.295 ;
        RECT 5.330 72.025 1204.470 74.855 ;
        RECT 5.330 66.585 1204.470 69.415 ;
        RECT 5.330 61.145 1204.470 63.975 ;
        RECT 5.330 55.705 1204.470 58.535 ;
        RECT 5.330 50.265 1204.470 53.095 ;
        RECT 5.330 44.825 1204.470 47.655 ;
        RECT 5.330 39.385 1204.470 42.215 ;
        RECT 5.330 33.945 1204.470 36.775 ;
        RECT 5.330 28.505 1204.470 31.335 ;
        RECT 5.330 23.065 1204.470 25.895 ;
        RECT 5.330 17.625 1204.470 20.455 ;
        RECT 5.330 12.185 1204.470 15.015 ;
      LAYER li1 ;
        RECT 5.520 10.795 1204.280 1498.805 ;
      LAYER met1 ;
        RECT 5.520 10.640 1204.280 1498.960 ;
      LAYER met2 ;
        RECT 21.070 1505.720 150.690 1506.610 ;
        RECT 151.530 1505.720 452.910 1506.610 ;
        RECT 453.750 1505.720 755.590 1506.610 ;
        RECT 756.430 1505.720 1057.810 1506.610 ;
        RECT 1058.650 1505.720 1200.970 1506.610 ;
        RECT 21.070 4.280 1200.970 1505.720 ;
        RECT 21.070 3.670 150.690 4.280 ;
        RECT 151.530 3.670 452.910 4.280 ;
        RECT 453.750 3.670 755.590 4.280 ;
        RECT 756.430 3.670 1057.810 4.280 ;
        RECT 1058.650 3.670 1200.970 4.280 ;
      LAYER met3 ;
        RECT 21.040 755.840 1206.000 1498.885 ;
        RECT 21.040 754.440 1205.600 755.840 ;
        RECT 21.040 10.715 1206.000 754.440 ;
      LAYER met4 ;
        RECT 637.855 537.375 711.840 952.505 ;
        RECT 714.240 537.375 788.640 952.505 ;
        RECT 791.040 537.375 865.440 952.505 ;
        RECT 867.840 537.375 930.745 952.505 ;
  END
END grp_99_SPI_TapeOutBlockRTL_32bits_5entries
END LIBRARY


magic
tech sky130A
magscale 1 2
timestamp 1655481716
<< obsli1 >>
rect 1104 2159 178848 177361
<< obsm1 >>
rect 1104 2128 178848 177392
<< metal2 >>
rect 15014 179200 15070 180000
rect 45006 179200 45062 180000
rect 74998 179200 75054 180000
rect 104990 179200 105046 180000
rect 134982 179200 135038 180000
rect 164974 179200 165030 180000
rect 17958 0 18014 800
rect 53930 0 53986 800
rect 89902 0 89958 800
rect 125966 0 126022 800
rect 161938 0 161994 800
<< obsm2 >>
rect 1398 179144 14958 179330
rect 15126 179144 44950 179330
rect 45118 179144 74942 179330
rect 75110 179144 104934 179330
rect 105102 179144 134926 179330
rect 135094 179144 164918 179330
rect 165086 179144 178186 179330
rect 1398 856 178186 179144
rect 1398 800 17902 856
rect 18070 800 53874 856
rect 54042 800 89846 856
rect 90014 800 125910 856
rect 126078 800 161882 856
rect 162050 800 178186 856
<< metal3 >>
rect 0 157496 800 157616
rect 179200 149880 180000 150000
rect 0 112480 800 112600
rect 179200 89904 180000 90024
rect 0 67464 800 67584
rect 179200 29928 180000 30048
rect 0 22448 800 22568
<< obsm3 >>
rect 800 157696 179200 177377
rect 880 157416 179200 157696
rect 800 150080 179200 157416
rect 800 149800 179120 150080
rect 800 112680 179200 149800
rect 880 112400 179200 112680
rect 800 90104 179200 112400
rect 800 89824 179120 90104
rect 800 67664 179200 89824
rect 880 67384 179200 67664
rect 800 30128 179200 67384
rect 800 29848 179120 30128
rect 800 22648 179200 29848
rect 880 22368 179200 22648
rect 800 2143 179200 22368
<< metal4 >>
rect 4208 2128 4528 177392
rect 19568 2128 19888 177392
rect 34928 2128 35248 177392
rect 50288 2128 50608 177392
rect 65648 2128 65968 177392
rect 81008 2128 81328 177392
rect 96368 2128 96688 177392
rect 111728 2128 112048 177392
rect 127088 2128 127408 177392
rect 142448 2128 142768 177392
rect 157808 2128 158128 177392
rect 173168 2128 173488 177392
<< labels >>
rlabel metal2 s 89902 0 89958 800 6 adapter_parity
port 1 nsew signal output
rlabel metal2 s 134982 179200 135038 180000 6 ap_en
port 2 nsew signal output
rlabel metal2 s 15014 179200 15070 180000 6 clk
port 3 nsew signal input
rlabel metal2 s 45006 179200 45062 180000 6 clk_en
port 4 nsew signal output
rlabel metal2 s 164974 179200 165030 180000 6 cs_en
port 5 nsew signal output
rlabel metal2 s 17958 0 18014 800 6 loopthrough_sel
port 6 nsew signal input
rlabel metal3 s 0 112480 800 112600 6 lt_sel_en
port 7 nsew signal output
rlabel metal2 s 53930 0 53986 800 6 minion_parity
port 8 nsew signal output
rlabel metal3 s 0 157496 800 157616 6 miso_en
port 9 nsew signal output
rlabel metal3 s 179200 149880 180000 150000 6 mosi_en
port 10 nsew signal output
rlabel metal2 s 125966 0 126022 800 6 mp_en
port 11 nsew signal output
rlabel metal2 s 74998 179200 75054 180000 6 reset
port 12 nsew signal input
rlabel metal2 s 104990 179200 105046 180000 6 reset_en
port 13 nsew signal output
rlabel metal2 s 161938 0 161994 800 6 sclk_en
port 14 nsew signal output
rlabel metal3 s 179200 29928 180000 30048 6 spi_min_cs
port 15 nsew signal input
rlabel metal3 s 0 67464 800 67584 6 spi_min_miso
port 16 nsew signal output
rlabel metal3 s 0 22448 800 22568 6 spi_min_mosi
port 17 nsew signal input
rlabel metal3 s 179200 89904 180000 90024 6 spi_min_sclk
port 18 nsew signal input
rlabel metal4 s 4208 2128 4528 177392 6 vccd1
port 19 nsew power input
rlabel metal4 s 34928 2128 35248 177392 6 vccd1
port 19 nsew power input
rlabel metal4 s 65648 2128 65968 177392 6 vccd1
port 19 nsew power input
rlabel metal4 s 96368 2128 96688 177392 6 vccd1
port 19 nsew power input
rlabel metal4 s 127088 2128 127408 177392 6 vccd1
port 19 nsew power input
rlabel metal4 s 157808 2128 158128 177392 6 vccd1
port 19 nsew power input
rlabel metal4 s 19568 2128 19888 177392 6 vssd1
port 20 nsew ground input
rlabel metal4 s 50288 2128 50608 177392 6 vssd1
port 20 nsew ground input
rlabel metal4 s 81008 2128 81328 177392 6 vssd1
port 20 nsew ground input
rlabel metal4 s 111728 2128 112048 177392 6 vssd1
port 20 nsew ground input
rlabel metal4 s 142448 2128 142768 177392 6 vssd1
port 20 nsew ground input
rlabel metal4 s 173168 2128 173488 177392 6 vssd1
port 20 nsew ground input
<< properties >>
string FIXED_BBOX 0 0 180000 180000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 16087492
string GDS_FILE /home/acm289/ece5745-tapeout/openlane/project-group15/runs/project-group15/results/finishing/grp_15_SPI_TapeOutBlockRTL_32bits_5entries.magic.gds
string GDS_START 641972
<< end >>


magic
tech sky130A
magscale 1 2
timestamp 1654279947
<< obsli1 >>
rect 1104 2159 240856 299761
<< obsm1 >>
rect 1104 2128 240856 299792
<< metal2 >>
rect 30194 301200 30250 302000
rect 90638 301200 90694 302000
rect 151174 301200 151230 302000
rect 211618 301200 211674 302000
rect 24214 0 24270 800
rect 72606 0 72662 800
rect 120998 0 121054 800
rect 169390 0 169446 800
rect 217782 0 217838 800
<< obsm2 >>
rect 1398 301144 30138 301322
rect 30306 301144 90582 301322
rect 90750 301144 151118 301322
rect 151286 301144 211562 301322
rect 211730 301144 240194 301322
rect 1398 856 240194 301144
rect 1398 800 24158 856
rect 24326 800 72550 856
rect 72718 800 120942 856
rect 121110 800 169334 856
rect 169502 800 217726 856
rect 217894 800 240194 856
<< metal3 >>
rect 241200 280304 242000 280424
rect 241200 237192 242000 237312
rect 0 226448 800 226568
rect 241200 194080 242000 194200
rect 241200 150832 242000 150952
rect 241200 107720 242000 107840
rect 0 75488 800 75608
rect 241200 64608 242000 64728
rect 241200 21496 242000 21616
<< obsm3 >>
rect 800 280504 241200 299777
rect 800 280224 241120 280504
rect 800 237392 241200 280224
rect 800 237112 241120 237392
rect 800 226648 241200 237112
rect 880 226368 241200 226648
rect 800 194280 241200 226368
rect 800 194000 241120 194280
rect 800 151032 241200 194000
rect 800 150752 241120 151032
rect 800 107920 241200 150752
rect 800 107640 241120 107920
rect 800 75688 241200 107640
rect 880 75408 241200 75688
rect 800 64808 241200 75408
rect 800 64528 241120 64808
rect 800 21696 241200 64528
rect 800 21416 241120 21696
rect 800 2143 241200 21416
<< metal4 >>
rect 4208 2128 4528 299792
rect 19568 2128 19888 299792
rect 34928 2128 35248 299792
rect 50288 2128 50608 299792
rect 65648 2128 65968 299792
rect 81008 2128 81328 299792
rect 96368 2128 96688 299792
rect 111728 2128 112048 299792
rect 127088 2128 127408 299792
rect 142448 2128 142768 299792
rect 157808 2128 158128 299792
rect 173168 2128 173488 299792
rect 188528 2128 188848 299792
rect 203888 2128 204208 299792
rect 219248 2128 219568 299792
rect 234608 2128 234928 299792
<< obsm4 >>
rect 113403 191251 127008 254285
rect 127488 191251 142368 254285
rect 142848 191251 157728 254285
rect 158208 191251 173088 254285
rect 173568 191251 179893 254285
<< labels >>
rlabel metal2 s 151174 301200 151230 302000 6 adapter_parity
port 1 nsew signal output
rlabel metal3 s 241200 194080 242000 194200 6 ap_en
port 2 nsew signal output
rlabel metal2 s 24214 0 24270 800 6 clk
port 3 nsew signal input
rlabel metal2 s 72606 0 72662 800 6 clk_en
port 4 nsew signal output
rlabel metal3 s 241200 21496 242000 21616 6 cs_en
port 5 nsew signal output
rlabel metal2 s 30194 301200 30250 302000 6 loopthrough_sel
port 6 nsew signal input
rlabel metal2 s 217782 0 217838 800 6 lt_sel_en
port 7 nsew signal output
rlabel metal2 s 90638 301200 90694 302000 6 minion_parity
port 8 nsew signal output
rlabel metal3 s 241200 64608 242000 64728 6 miso_en
port 9 nsew signal output
rlabel metal3 s 241200 107720 242000 107840 6 mosi_en
port 10 nsew signal output
rlabel metal3 s 0 75488 800 75608 6 mp_en
port 11 nsew signal output
rlabel metal2 s 120998 0 121054 800 6 reset
port 12 nsew signal input
rlabel metal2 s 169390 0 169446 800 6 reset_en
port 13 nsew signal output
rlabel metal3 s 241200 150832 242000 150952 6 sclk_en
port 14 nsew signal output
rlabel metal2 s 211618 301200 211674 302000 6 spi_min__cs
port 15 nsew signal input
rlabel metal3 s 241200 237192 242000 237312 6 spi_min__miso
port 16 nsew signal output
rlabel metal3 s 0 226448 800 226568 6 spi_min__mosi
port 17 nsew signal input
rlabel metal3 s 241200 280304 242000 280424 6 spi_min__sclk
port 18 nsew signal input
rlabel metal4 s 4208 2128 4528 299792 6 vccd1
port 19 nsew power input
rlabel metal4 s 34928 2128 35248 299792 6 vccd1
port 19 nsew power input
rlabel metal4 s 65648 2128 65968 299792 6 vccd1
port 19 nsew power input
rlabel metal4 s 96368 2128 96688 299792 6 vccd1
port 19 nsew power input
rlabel metal4 s 127088 2128 127408 299792 6 vccd1
port 19 nsew power input
rlabel metal4 s 157808 2128 158128 299792 6 vccd1
port 19 nsew power input
rlabel metal4 s 188528 2128 188848 299792 6 vccd1
port 19 nsew power input
rlabel metal4 s 219248 2128 219568 299792 6 vccd1
port 19 nsew power input
rlabel metal4 s 19568 2128 19888 299792 6 vssd1
port 20 nsew ground input
rlabel metal4 s 50288 2128 50608 299792 6 vssd1
port 20 nsew ground input
rlabel metal4 s 81008 2128 81328 299792 6 vssd1
port 20 nsew ground input
rlabel metal4 s 111728 2128 112048 299792 6 vssd1
port 20 nsew ground input
rlabel metal4 s 142448 2128 142768 299792 6 vssd1
port 20 nsew ground input
rlabel metal4 s 173168 2128 173488 299792 6 vssd1
port 20 nsew ground input
rlabel metal4 s 203888 2128 204208 299792 6 vssd1
port 20 nsew ground input
rlabel metal4 s 234608 2128 234928 299792 6 vssd1
port 20 nsew ground input
<< properties >>
string FIXED_BBOX 0 0 242000 302000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 27708114
string GDS_FILE /home/acm289/ece5745-tapeout/openlane/project-group99/runs/project-group99/results/finishing/grp_99_SPI_TapeOutBlockRTL_32bits_5entries.magic.gds
string GDS_START 472510
<< end >>


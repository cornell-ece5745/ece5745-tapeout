magic
tech sky130A
magscale 1 2
timestamp 1654706468
<< obsli1 >>
rect 1104 2159 240856 299761
<< obsm1 >>
rect 1104 2128 240856 299792
<< metal2 >>
rect 40314 301200 40370 302000
rect 120906 301200 120962 302000
rect 201590 301200 201646 302000
rect 15106 0 15162 800
rect 45282 0 45338 800
rect 75550 0 75606 800
rect 105818 0 105874 800
rect 136086 0 136142 800
rect 166262 0 166318 800
rect 196530 0 196586 800
rect 226798 0 226854 800
<< obsm2 >>
rect 1398 301144 40258 301322
rect 40426 301144 120850 301322
rect 121018 301144 201534 301322
rect 201702 301144 240194 301322
rect 1398 856 240194 301144
rect 1398 800 15050 856
rect 15218 800 45226 856
rect 45394 800 75494 856
rect 75662 800 105762 856
rect 105930 800 136030 856
rect 136198 800 166206 856
rect 166374 800 196474 856
rect 196642 800 226742 856
rect 226910 800 240194 856
<< metal3 >>
rect 241200 271736 242000 271856
rect 0 226448 800 226568
rect 241200 211352 242000 211472
rect 241200 150968 242000 151088
rect 241200 90584 242000 90704
rect 0 75488 800 75608
rect 241200 30200 242000 30320
<< obsm3 >>
rect 800 271936 241200 299777
rect 800 271656 241120 271936
rect 800 226648 241200 271656
rect 880 226368 241200 226648
rect 800 211552 241200 226368
rect 800 211272 241120 211552
rect 800 151168 241200 211272
rect 800 150888 241120 151168
rect 800 90784 241200 150888
rect 800 90504 241120 90784
rect 800 75688 241200 90504
rect 880 75408 241200 75688
rect 800 30400 241200 75408
rect 800 30120 241120 30400
rect 800 2143 241200 30120
<< metal4 >>
rect 4208 2128 4528 299792
rect 19568 2128 19888 299792
rect 34928 2128 35248 299792
rect 50288 2128 50608 299792
rect 65648 2128 65968 299792
rect 81008 2128 81328 299792
rect 96368 2128 96688 299792
rect 111728 2128 112048 299792
rect 127088 2128 127408 299792
rect 142448 2128 142768 299792
rect 157808 2128 158128 299792
rect 173168 2128 173488 299792
rect 188528 2128 188848 299792
rect 203888 2128 204208 299792
rect 219248 2128 219568 299792
rect 234608 2128 234928 299792
<< obsm4 >>
rect 138427 3435 142368 176901
rect 142848 3435 157728 176901
rect 158208 3435 173088 176901
rect 173568 3435 188448 176901
rect 188928 3435 193141 176901
<< labels >>
rlabel metal2 s 201590 301200 201646 302000 6 adapter_parity
port 1 nsew signal output
rlabel metal2 s 136086 0 136142 800 6 ap_en
port 2 nsew signal output
rlabel metal2 s 15106 0 15162 800 6 clk
port 3 nsew signal input
rlabel metal2 s 45282 0 45338 800 6 clk_en
port 4 nsew signal output
rlabel metal3 s 241200 30200 242000 30320 6 cs_en
port 5 nsew signal output
rlabel metal2 s 40314 301200 40370 302000 6 loopthrough_sel
port 6 nsew signal input
rlabel metal3 s 0 75488 800 75608 6 lt_sel_en
port 7 nsew signal output
rlabel metal2 s 120906 301200 120962 302000 6 minion_parity
port 8 nsew signal output
rlabel metal3 s 241200 90584 242000 90704 6 miso_en
port 9 nsew signal output
rlabel metal3 s 241200 150968 242000 151088 6 mosi_en
port 10 nsew signal output
rlabel metal3 s 0 226448 800 226568 6 mp_en
port 11 nsew signal output
rlabel metal2 s 75550 0 75606 800 6 reset
port 12 nsew signal input
rlabel metal2 s 105818 0 105874 800 6 reset_en
port 13 nsew signal output
rlabel metal3 s 241200 211352 242000 211472 6 sclk_en
port 14 nsew signal output
rlabel metal2 s 166262 0 166318 800 6 spi_min__cs
port 15 nsew signal input
rlabel metal2 s 196530 0 196586 800 6 spi_min__miso
port 16 nsew signal output
rlabel metal3 s 241200 271736 242000 271856 6 spi_min__mosi
port 17 nsew signal input
rlabel metal2 s 226798 0 226854 800 6 spi_min__sclk
port 18 nsew signal input
rlabel metal4 s 4208 2128 4528 299792 6 vccd1
port 19 nsew power input
rlabel metal4 s 34928 2128 35248 299792 6 vccd1
port 19 nsew power input
rlabel metal4 s 65648 2128 65968 299792 6 vccd1
port 19 nsew power input
rlabel metal4 s 96368 2128 96688 299792 6 vccd1
port 19 nsew power input
rlabel metal4 s 127088 2128 127408 299792 6 vccd1
port 19 nsew power input
rlabel metal4 s 157808 2128 158128 299792 6 vccd1
port 19 nsew power input
rlabel metal4 s 188528 2128 188848 299792 6 vccd1
port 19 nsew power input
rlabel metal4 s 219248 2128 219568 299792 6 vccd1
port 19 nsew power input
rlabel metal4 s 19568 2128 19888 299792 6 vssd1
port 20 nsew ground input
rlabel metal4 s 50288 2128 50608 299792 6 vssd1
port 20 nsew ground input
rlabel metal4 s 81008 2128 81328 299792 6 vssd1
port 20 nsew ground input
rlabel metal4 s 111728 2128 112048 299792 6 vssd1
port 20 nsew ground input
rlabel metal4 s 142448 2128 142768 299792 6 vssd1
port 20 nsew ground input
rlabel metal4 s 173168 2128 173488 299792 6 vssd1
port 20 nsew ground input
rlabel metal4 s 203888 2128 204208 299792 6 vssd1
port 20 nsew ground input
rlabel metal4 s 234608 2128 234928 299792 6 vssd1
port 20 nsew ground input
<< properties >>
string FIXED_BBOX 0 0 242000 302000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 27341118
string GDS_FILE /home/acm289/ece5745-tapeout/openlane/project-group99/runs/project-group99/results/finishing/grp_99_SPI_TapeOutBlockRTL_32bits_5entries.magic.gds
string GDS_START 507378
<< end >>


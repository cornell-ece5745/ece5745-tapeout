VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO grp_99_SPI_TapeOutBlockRTL_32bits_5entries
  CLASS BLOCK ;
  FOREIGN grp_99_SPI_TapeOutBlockRTL_32bits_5entries ;
  ORIGIN 0.000 0.000 ;
  SIZE 1210.000 BY 1510.000 ;
  PIN adapter_parity
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1007.950 1506.000 1008.230 1510.000 ;
    END
  END adapter_parity
  PIN ap_en
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 680.430 0.000 680.710 4.000 ;
    END
  END ap_en
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.530 0.000 75.810 4.000 ;
    END
  END clk
  PIN clk_en
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 226.410 0.000 226.690 4.000 ;
    END
  END clk_en
  PIN cs_en
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1206.000 151.000 1210.000 151.600 ;
    END
  END cs_en
  PIN loopthrough_sel
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 201.570 1506.000 201.850 1510.000 ;
    END
  END loopthrough_sel
  PIN lt_sel_en
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 377.440 4.000 378.040 ;
    END
  END lt_sel_en
  PIN minion_parity
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 604.530 1506.000 604.810 1510.000 ;
    END
  END minion_parity
  PIN miso_en
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1206.000 452.920 1210.000 453.520 ;
    END
  END miso_en
  PIN mosi_en
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1206.000 754.840 1210.000 755.440 ;
    END
  END mosi_en
  PIN mp_en
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1132.240 4.000 1132.840 ;
    END
  END mp_en
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 377.750 0.000 378.030 4.000 ;
    END
  END reset
  PIN reset_en
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 529.090 0.000 529.370 4.000 ;
    END
  END reset_en
  PIN sclk_en
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1206.000 1056.760 1210.000 1057.360 ;
    END
  END sclk_en
  PIN spi_min__cs
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 831.310 0.000 831.590 4.000 ;
    END
  END spi_min__cs
  PIN spi_min__miso
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 982.650 0.000 982.930 4.000 ;
    END
  END spi_min__miso
  PIN spi_min__mosi
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1206.000 1358.680 1210.000 1359.280 ;
    END
  END spi_min__mosi
  PIN spi_min__sclk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1133.990 0.000 1134.270 4.000 ;
    END
  END spi_min__sclk
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 1498.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 1498.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 1498.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 1498.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 1498.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 1498.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 942.640 10.640 944.240 1498.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 1096.240 10.640 1097.840 1498.960 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 1498.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 1498.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 1498.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 1498.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 1498.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 1498.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 1019.440 10.640 1021.040 1498.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 1173.040 10.640 1174.640 1498.960 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 1204.280 1498.805 ;
      LAYER met1 ;
        RECT 5.520 10.640 1204.280 1498.960 ;
      LAYER met2 ;
        RECT 6.990 1505.720 201.290 1506.610 ;
        RECT 202.130 1505.720 604.250 1506.610 ;
        RECT 605.090 1505.720 1007.670 1506.610 ;
        RECT 1008.510 1505.720 1200.970 1506.610 ;
        RECT 6.990 4.280 1200.970 1505.720 ;
        RECT 6.990 4.000 75.250 4.280 ;
        RECT 76.090 4.000 226.130 4.280 ;
        RECT 226.970 4.000 377.470 4.280 ;
        RECT 378.310 4.000 528.810 4.280 ;
        RECT 529.650 4.000 680.150 4.280 ;
        RECT 680.990 4.000 831.030 4.280 ;
        RECT 831.870 4.000 982.370 4.280 ;
        RECT 983.210 4.000 1133.710 4.280 ;
        RECT 1134.550 4.000 1200.970 4.280 ;
      LAYER met3 ;
        RECT 4.000 1359.680 1206.000 1498.885 ;
        RECT 4.000 1358.280 1205.600 1359.680 ;
        RECT 4.000 1133.240 1206.000 1358.280 ;
        RECT 4.400 1131.840 1206.000 1133.240 ;
        RECT 4.000 1057.760 1206.000 1131.840 ;
        RECT 4.000 1056.360 1205.600 1057.760 ;
        RECT 4.000 755.840 1206.000 1056.360 ;
        RECT 4.000 754.440 1205.600 755.840 ;
        RECT 4.000 453.920 1206.000 754.440 ;
        RECT 4.000 452.520 1205.600 453.920 ;
        RECT 4.000 378.440 1206.000 452.520 ;
        RECT 4.400 377.040 1206.000 378.440 ;
        RECT 4.000 152.000 1206.000 377.040 ;
        RECT 4.000 150.600 1205.600 152.000 ;
        RECT 4.000 10.715 1206.000 150.600 ;
      LAYER met4 ;
        RECT 692.135 17.175 711.840 884.505 ;
        RECT 714.240 17.175 788.640 884.505 ;
        RECT 791.040 17.175 865.440 884.505 ;
        RECT 867.840 17.175 942.240 884.505 ;
        RECT 944.640 17.175 965.705 884.505 ;
  END
END grp_99_SPI_TapeOutBlockRTL_32bits_5entries
END LIBRARY


magic
tech sky130A
magscale 1 2
timestamp 1655317030
<< obsli1 >>
rect 1104 2159 240856 299761
<< obsm1 >>
rect 1104 2128 240856 299792
<< metal2 >>
rect 40314 301200 40370 302000
rect 120906 301200 120962 302000
rect 201590 301200 201646 302000
rect 20166 0 20222 800
rect 60462 0 60518 800
rect 100758 0 100814 800
rect 141146 0 141202 800
rect 181442 0 181498 800
rect 221738 0 221794 800
<< obsm2 >>
rect 1398 301144 40258 301322
rect 40426 301144 120850 301322
rect 121018 301144 201534 301322
rect 201702 301144 240194 301322
rect 1398 856 240194 301144
rect 1398 734 20110 856
rect 20278 734 60406 856
rect 60574 734 100702 856
rect 100870 734 141090 856
rect 141258 734 181386 856
rect 181554 734 221682 856
rect 221850 734 240194 856
<< metal3 >>
rect 241200 276768 242000 276888
rect 0 251608 800 251728
rect 241200 226448 242000 226568
rect 241200 176128 242000 176248
rect 0 150968 800 151088
rect 241200 125808 242000 125928
rect 241200 75488 242000 75608
rect 0 50328 800 50448
rect 241200 25168 242000 25288
<< obsm3 >>
rect 800 276968 241200 299777
rect 800 276688 241120 276968
rect 800 251808 241200 276688
rect 880 251528 241200 251808
rect 800 226648 241200 251528
rect 800 226368 241120 226648
rect 800 176328 241200 226368
rect 800 176048 241120 176328
rect 800 151168 241200 176048
rect 880 150888 241200 151168
rect 800 126008 241200 150888
rect 800 125728 241120 126008
rect 800 75688 241200 125728
rect 800 75408 241120 75688
rect 800 50528 241200 75408
rect 880 50248 241200 50528
rect 800 25368 241200 50248
rect 800 25088 241120 25368
rect 800 2143 241200 25088
<< metal4 >>
rect 4208 2128 4528 299792
rect 19568 2128 19888 299792
rect 34928 2128 35248 299792
rect 50288 2128 50608 299792
rect 65648 2128 65968 299792
rect 81008 2128 81328 299792
rect 96368 2128 96688 299792
rect 111728 2128 112048 299792
rect 127088 2128 127408 299792
rect 142448 2128 142768 299792
rect 157808 2128 158128 299792
rect 173168 2128 173488 299792
rect 188528 2128 188848 299792
rect 203888 2128 204208 299792
rect 219248 2128 219568 299792
rect 234608 2128 234928 299792
<< obsm4 >>
rect 102179 140659 111648 233749
rect 112128 140659 127008 233749
rect 127488 140659 142368 233749
rect 142848 140659 157728 233749
rect 158208 140659 173088 233749
rect 173568 140659 175845 233749
<< labels >>
rlabel metal2 s 201590 301200 201646 302000 6 adapter_parity
port 1 nsew signal output
rlabel metal2 s 181442 0 181498 800 6 ap_en
port 2 nsew signal output
rlabel metal2 s 20166 0 20222 800 6 clk
port 3 nsew signal input
rlabel metal2 s 60462 0 60518 800 6 clk_en
port 4 nsew signal output
rlabel metal3 s 241200 25168 242000 25288 6 cs_en
port 5 nsew signal output
rlabel metal2 s 40314 301200 40370 302000 6 loopthrough_sel
port 6 nsew signal input
rlabel metal3 s 0 50328 800 50448 6 lt_sel_en
port 7 nsew signal output
rlabel metal2 s 120906 301200 120962 302000 6 minion_parity
port 8 nsew signal output
rlabel metal3 s 241200 75488 242000 75608 6 miso_en
port 9 nsew signal output
rlabel metal3 s 241200 125808 242000 125928 6 mosi_en
port 10 nsew signal output
rlabel metal3 s 0 150968 800 151088 6 mp_en
port 11 nsew signal output
rlabel metal2 s 100758 0 100814 800 6 reset
port 12 nsew signal input
rlabel metal2 s 141146 0 141202 800 6 reset_en
port 13 nsew signal output
rlabel metal3 s 241200 176128 242000 176248 6 sclk_en
port 14 nsew signal output
rlabel metal3 s 241200 226448 242000 226568 6 spi_min__cs
port 15 nsew signal input
rlabel metal2 s 221738 0 221794 800 6 spi_min__miso
port 16 nsew signal output
rlabel metal3 s 0 251608 800 251728 6 spi_min__mosi
port 17 nsew signal input
rlabel metal3 s 241200 276768 242000 276888 6 spi_min__sclk
port 18 nsew signal input
rlabel metal4 s 4208 2128 4528 299792 6 vccd1
port 19 nsew power input
rlabel metal4 s 34928 2128 35248 299792 6 vccd1
port 19 nsew power input
rlabel metal4 s 65648 2128 65968 299792 6 vccd1
port 19 nsew power input
rlabel metal4 s 96368 2128 96688 299792 6 vccd1
port 19 nsew power input
rlabel metal4 s 127088 2128 127408 299792 6 vccd1
port 19 nsew power input
rlabel metal4 s 157808 2128 158128 299792 6 vccd1
port 19 nsew power input
rlabel metal4 s 188528 2128 188848 299792 6 vccd1
port 19 nsew power input
rlabel metal4 s 219248 2128 219568 299792 6 vccd1
port 19 nsew power input
rlabel metal4 s 19568 2128 19888 299792 6 vssd1
port 20 nsew ground input
rlabel metal4 s 50288 2128 50608 299792 6 vssd1
port 20 nsew ground input
rlabel metal4 s 81008 2128 81328 299792 6 vssd1
port 20 nsew ground input
rlabel metal4 s 111728 2128 112048 299792 6 vssd1
port 20 nsew ground input
rlabel metal4 s 142448 2128 142768 299792 6 vssd1
port 20 nsew ground input
rlabel metal4 s 173168 2128 173488 299792 6 vssd1
port 20 nsew ground input
rlabel metal4 s 203888 2128 204208 299792 6 vssd1
port 20 nsew ground input
rlabel metal4 s 234608 2128 234928 299792 6 vssd1
port 20 nsew ground input
<< properties >>
string FIXED_BBOX 0 0 242000 302000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 29895272
string GDS_FILE /home/acm289/ece5745-tapeout/openlane/project-group99/runs/project-group99/results/finishing/grp_99_SPI_TapeOutBlockRTL_32bits_5entries.magic.gds
string GDS_START 661568
<< end >>


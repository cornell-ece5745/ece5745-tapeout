
//------> /opt/MentorGraphics/catapult/pkgs/siflibs/ccs_in_wait_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module ccs_in_wait_v1 (idat, rdy, ivld, dat, irdy, vld);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  output             rdy;
  output             ivld;
  input  [width-1:0] dat;
  input              irdy;
  input              vld;

  wire   [width-1:0] idat;
  wire               rdy;
  wire               ivld;

  localparam stallOff = 0; 
  wire                  stall_ctrl;
  assign stall_ctrl = stallOff;

  assign idat = dat;
  assign rdy = irdy && !stall_ctrl;
  assign ivld = vld && !stall_ctrl;

endmodule


//------> /opt/MentorGraphics/catapult/pkgs/siflibs/ccs_out_wait_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module ccs_out_wait_v1 (dat, irdy, vld, idat, rdy, ivld);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] dat;
  output             irdy;
  output             vld;
  input  [width-1:0] idat;
  input              rdy;
  input              ivld;

  wire   [width-1:0] dat;
  wire               irdy;
  wire               vld;

  localparam stallOff = 0; 
  wire stall_ctrl;
  assign stall_ctrl = stallOff;

  assign dat = idat;
  assign irdy = rdy && !stall_ctrl;
  assign vld = ivld && !stall_ctrl;

endmodule



//------> ./rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    2021.1/950854 Production Release
//  HLS Date:       Mon Aug  2 21:36:02 PDT 2021
// 
//  Generated by:   tdt46@en-ec-ecelinux-01.coecis.cornell.edu
//  Generated date: Sat May 21 19:05:18 2022
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    crc32_core_core_fsm
//  FSM Module
// ------------------------------------------------------------------


module crc32_core_core_fsm (
  clk, rst, core_wen, fsm_output, main_C_0_tr0, for_C_0_tr0
);
  input clk;
  input rst;
  input core_wen;
  output [3:0] fsm_output;
  reg [3:0] fsm_output;
  input main_C_0_tr0;
  input for_C_0_tr0;


  // FSM State Type Declaration for crc32_core_core_fsm_1
  parameter
    core_rlp_C_0 = 2'd0,
    main_C_0 = 2'd1,
    for_C_0 = 2'd2,
    main_C_1 = 2'd3;

  reg [1:0] state_var;
  reg [1:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : crc32_core_core_fsm_1
    case (state_var)
      main_C_0 : begin
        fsm_output = 4'b0010;
        if ( main_C_0_tr0 ) begin
          state_var_NS = main_C_1;
        end
        else begin
          state_var_NS = for_C_0;
        end
      end
      for_C_0 : begin
        fsm_output = 4'b0100;
        if ( for_C_0_tr0 ) begin
          state_var_NS = main_C_1;
        end
        else begin
          state_var_NS = for_C_0;
        end
      end
      main_C_1 : begin
        fsm_output = 4'b1000;
        state_var_NS = main_C_0;
      end
      // core_rlp_C_0
      default : begin
        fsm_output = 4'b0001;
        state_var_NS = main_C_0;
      end
    endcase
  end

  always @(posedge clk) begin
    if ( rst ) begin
      state_var <= core_rlp_C_0;
    end
    else if ( core_wen ) begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    crc32_core_staller
// ------------------------------------------------------------------


module crc32_core_staller (
  core_wen, in_rsci_wen_comp, out_rsci_wen_comp
);
  output core_wen;
  input in_rsci_wen_comp;
  input out_rsci_wen_comp;



  // Interconnect Declarations for Component Instantiations 
  assign core_wen = in_rsci_wen_comp & out_rsci_wen_comp;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    crc32_core_out_rsci_out_wait_ctrl
// ------------------------------------------------------------------


module crc32_core_out_rsci_out_wait_ctrl (
  out_rsci_iswt0, out_rsci_biwt, out_rsci_irdy
);
  input out_rsci_iswt0;
  output out_rsci_biwt;
  input out_rsci_irdy;



  // Interconnect Declarations for Component Instantiations 
  assign out_rsci_biwt = out_rsci_iswt0 & out_rsci_irdy;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    crc32_core_in_rsci_in_wait_ctrl
// ------------------------------------------------------------------


module crc32_core_in_rsci_in_wait_ctrl (
  in_rsci_iswt0, in_rsci_biwt, in_rsci_ivld
);
  input in_rsci_iswt0;
  output in_rsci_biwt;
  input in_rsci_ivld;



  // Interconnect Declarations for Component Instantiations 
  assign in_rsci_biwt = in_rsci_iswt0 & in_rsci_ivld;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    crc32_core_out_rsci
// ------------------------------------------------------------------


module crc32_core_out_rsci (
  out_rsc_dat, out_rsc_vld, out_rsc_rdy, out_rsci_oswt, out_rsci_wen_comp, out_rsci_idat
);
  output [31:0] out_rsc_dat;
  output out_rsc_vld;
  input out_rsc_rdy;
  input out_rsci_oswt;
  output out_rsci_wen_comp;
  input [31:0] out_rsci_idat;


  // Interconnect Declarations
  wire out_rsci_biwt;
  wire out_rsci_irdy;


  // Interconnect Declarations for Component Instantiations 
  ccs_out_wait_v1 #(.rscid(32'sd2),
  .width(32'sd32)) out_rsci (
      .irdy(out_rsci_irdy),
      .ivld(out_rsci_oswt),
      .idat(out_rsci_idat),
      .rdy(out_rsc_rdy),
      .vld(out_rsc_vld),
      .dat(out_rsc_dat)
    );
  crc32_core_out_rsci_out_wait_ctrl crc32_core_out_rsci_out_wait_ctrl_inst (
      .out_rsci_iswt0(out_rsci_oswt),
      .out_rsci_biwt(out_rsci_biwt),
      .out_rsci_irdy(out_rsci_irdy)
    );
  assign out_rsci_wen_comp = (~ out_rsci_oswt) | out_rsci_biwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    crc32_core_in_rsci
// ------------------------------------------------------------------


module crc32_core_in_rsci (
  in_rsc_dat, in_rsc_vld, in_rsc_rdy, in_rsci_oswt, in_rsci_wen_comp, in_rsci_idat_mxwt
);
  input [7:0] in_rsc_dat;
  input in_rsc_vld;
  output in_rsc_rdy;
  input in_rsci_oswt;
  output in_rsci_wen_comp;
  output [7:0] in_rsci_idat_mxwt;


  // Interconnect Declarations
  wire in_rsci_biwt;
  wire in_rsci_ivld;
  wire [7:0] in_rsci_idat;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_wait_v1 #(.rscid(32'sd1),
  .width(32'sd8)) in_rsci (
      .rdy(in_rsc_rdy),
      .vld(in_rsc_vld),
      .dat(in_rsc_dat),
      .irdy(in_rsci_oswt),
      .ivld(in_rsci_ivld),
      .idat(in_rsci_idat)
    );
  crc32_core_in_rsci_in_wait_ctrl crc32_core_in_rsci_in_wait_ctrl_inst (
      .in_rsci_iswt0(in_rsci_oswt),
      .in_rsci_biwt(in_rsci_biwt),
      .in_rsci_ivld(in_rsci_ivld)
    );
  assign in_rsci_idat_mxwt = in_rsci_idat;
  assign in_rsci_wen_comp = (~ in_rsci_oswt) | in_rsci_biwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    crc32_core
// ------------------------------------------------------------------


module crc32_core (
  clk, rst, in_rsc_dat, in_rsc_vld, in_rsc_rdy, out_rsc_dat, out_rsc_vld, out_rsc_rdy
);
  input clk;
  input rst;
  input [7:0] in_rsc_dat;
  input in_rsc_vld;
  output in_rsc_rdy;
  output [31:0] out_rsc_dat;
  output out_rsc_vld;
  input out_rsc_rdy;


  // Interconnect Declarations
  wire core_wen;
  wire in_rsci_wen_comp;
  wire [7:0] in_rsci_idat_mxwt;
  wire out_rsci_wen_comp;
  reg out_rsci_idat_31;
  reg out_rsci_idat_30;
  reg out_rsci_idat_29;
  reg out_rsci_idat_28;
  reg out_rsci_idat_27;
  reg out_rsci_idat_26;
  reg out_rsci_idat_25;
  reg out_rsci_idat_24;
  reg out_rsci_idat_23;
  reg out_rsci_idat_22;
  reg out_rsci_idat_21;
  reg out_rsci_idat_20;
  reg out_rsci_idat_19;
  reg out_rsci_idat_18;
  reg out_rsci_idat_17;
  reg out_rsci_idat_16;
  reg out_rsci_idat_15;
  reg out_rsci_idat_14;
  reg out_rsci_idat_13;
  reg out_rsci_idat_12;
  reg out_rsci_idat_11;
  reg out_rsci_idat_10;
  reg out_rsci_idat_9;
  reg out_rsci_idat_8;
  reg out_rsci_idat_7;
  reg out_rsci_idat_6;
  reg out_rsci_idat_5;
  reg out_rsci_idat_4;
  reg out_rsci_idat_3;
  reg out_rsci_idat_2;
  reg out_rsci_idat_1;
  reg out_rsci_idat_0;
  wire [3:0] fsm_output;
  wire for_for_8_b_xor_tmp;
  wire for_for_7_b_xor_tmp;
  wire for_for_6_b_xor_tmp;
  wire for_for_5_b_xor_tmp;
  wire for_for_4_b_xor_tmp;
  wire not_tmp_3;
  wire not_tmp_4;
  wire not_tmp_5;
  wire not_tmp_6;
  wire not_tmp_7;
  wire not_tmp_8;
  wire not_tmp_9;
  wire not_tmp_10;
  wire or_tmp_32;
  wire or_tmp_40;
  wire or_tmp_52;
  wire or_tmp_56;
  wire or_tmp_60;
  wire exit_for_sva_mx0;
  reg crc_2_1_sva;
  reg crc_1_1_sva;
  reg crc_0_1_sva;
  wire and_314_cse;
  reg reg_out_rsci_iswt0_cse;
  reg reg_in_rsci_iswt0_cse;
  wire crc_mux_140_cse;
  wire [8:0] z_out;
  wire [9:0] nl_z_out;
  reg [7:0] size_val_sva;
  reg crc_15_1_sva;
  reg crc_16_1_sva;
  reg crc_14_1_sva;
  reg crc_17_1_sva;
  reg crc_13_1_sva;
  reg crc_18_1_sva;
  reg crc_12_1_sva;
  reg crc_19_1_sva;
  reg crc_11_1_sva;
  reg crc_20_1_sva;
  reg crc_10_1_sva;
  reg crc_21_1_sva;
  reg crc_9_1_sva;
  reg crc_22_1_sva;
  reg crc_8_1_sva;
  reg crc_23_1_sva;
  reg crc_7_1_sva;
  reg crc_24_1_sva;
  reg crc_6_1_sva;
  reg crc_25_1_sva;
  reg crc_5_1_sva;
  reg crc_26_1_sva;
  reg crc_4_1_sva;
  reg crc_27_1_sva;
  reg crc_3_1_sva;
  reg crc_28_1_sva;
  reg crc_29_1_sva;
  reg crc_30_1_sva;
  reg crc_31_1_sva;
  reg [7:0] for_i_sva;
  wire crc_5_4_lpi_2_dfm_mx0;
  wire crc_8_2_lpi_2_dfm_mx0;
  wire crc_8_3_lpi_2_dfm_mx0;
  wire crc_8_4_lpi_2_dfm_mx0;
  wire crc_8_5_lpi_2_dfm_mx0;
  wire crc_8_6_lpi_2_dfm_mx0;
  wire crc_9_6_lpi_2_dfm_mx0;
  wire crc_9_7_lpi_2_dfm_mx0;
  wire crc_9_lpi_2_dfm_mx0;
  wire crc_15_3_lpi_2_dfm_mx0;
  wire crc_15_4_lpi_2_dfm_mx0;
  wire crc_15_5_lpi_2_dfm_mx0;
  wire crc_19_2_lpi_2_dfm_mx0;
  wire crc_19_3_lpi_2_dfm_mx0;
  wire crc_19_4_lpi_2_dfm_mx0;
  wire crc_19_5_lpi_2_dfm_mx0;
  wire crc_20_5_lpi_2_dfm_mx0;
  wire crc_20_6_lpi_2_dfm_mx0;
  wire crc_20_7_lpi_2_dfm_mx0;
  wire crc_20_lpi_2_dfm_mx0;
  wire crc_21_lpi_2_dfm_mx0;
  wire crc_23_7_lpi_2_dfm_mx0;
  wire crc_24_7_lpi_2_dfm_mx0;
  wire crc_24_lpi_2_dfm_mx0;
  wire crc_26_7_lpi_2_dfm_mx0;
  wire crc_27_7_lpi_2_dfm_mx0;
  wire crc_27_lpi_2_dfm_mx0;
  wire crc_29_7_lpi_2_dfm_mx0;
  wire crc_30_7_lpi_2_dfm_mx0;
  wire crc_30_lpi_2_dfm_mx0;
  wire for_for_b_2_sva_1;
  wire crc_15_2_lpi_2_dfm_mx0;
  wire crc_21_7_lpi_2_dfm_mx0;
  wire crc_23_6_lpi_2_dfm_mx0;
  wire crc_26_6_lpi_2_dfm_mx0;
  wire crc_29_6_lpi_2_dfm_mx0;
  wire for_for_b_1_sva_1;
  wire crc_21_6_lpi_2_dfm_mx0;
  wire crc_23_5_lpi_2_dfm_mx0;
  wire crc_24_6_lpi_2_dfm_mx0;
  wire crc_26_5_lpi_2_dfm_mx0;
  wire crc_27_6_lpi_2_dfm_mx0;
  wire crc_29_5_lpi_2_dfm_mx0;
  wire crc_30_6_lpi_2_dfm_mx0;
  wire crc_9_5_lpi_2_dfm_mx0;
  wire crc_21_5_lpi_2_dfm_mx0;
  wire crc_23_4_lpi_2_dfm_mx0;
  wire crc_24_5_lpi_2_dfm_mx0;
  wire crc_26_4_lpi_2_dfm_mx0;
  wire crc_27_5_lpi_2_dfm_mx0;
  wire crc_29_4_lpi_2_dfm_mx0;
  wire crc_30_5_lpi_2_dfm_mx0;
  wire crc_9_4_lpi_2_dfm_mx0;
  wire crc_20_4_lpi_2_dfm_mx0;
  wire crc_21_4_lpi_2_dfm_mx0;
  wire crc_23_3_lpi_2_dfm_mx0;
  wire crc_24_4_lpi_2_dfm_mx0;
  wire crc_26_3_lpi_2_dfm_mx0;
  wire crc_27_4_lpi_2_dfm_mx0;
  wire crc_29_3_lpi_2_dfm_mx0;
  wire crc_30_4_lpi_2_dfm_mx0;
  wire for_for_b_3_sva_1;
  wire crc_9_3_lpi_2_dfm_mx0;
  wire crc_20_3_lpi_2_dfm_mx0;
  wire crc_21_3_lpi_2_dfm_mx0;
  wire crc_23_2_lpi_2_dfm_mx0;
  wire crc_24_3_lpi_2_dfm_mx0;
  wire crc_26_2_lpi_2_dfm_mx0;
  wire crc_27_3_lpi_2_dfm_mx0;
  wire crc_29_2_lpi_2_dfm_mx0;
  wire crc_30_3_lpi_2_dfm_mx0;
  wire crc_9_2_lpi_2_dfm_mx0;
  wire crc_20_2_lpi_2_dfm_mx0;
  wire crc_21_2_lpi_2_dfm_mx0;
  wire crc_24_2_lpi_2_dfm_mx0;
  wire crc_27_2_lpi_2_dfm_mx0;
  wire crc_30_2_lpi_2_dfm_mx0;
  wire xor_cse_1;
  wire xor_cse_5;

  wire crc_mux_142_nl;
  wire crc_mux_144_nl;
  wire crc_mux_146_nl;
  wire crc_mux_148_nl;
  wire crc_mux_150_nl;
  wire crc_mux_152_nl;
  wire crc_mux_154_nl;
  wire crc_mux_156_nl;
  wire crc_mux_160_nl;
  wire crc_mux_162_nl;
  wire crc_mux_164_nl;
  wire crc_mux_166_nl;
  wire crc_mux_165_nl;
  wire crc_mux_163_nl;
  wire crc_mux_161_nl;
  wire crc_mux_159_nl;
  wire crc_mux_158_nl;
  wire crc_mux_157_nl;
  wire crc_mux_155_nl;
  wire crc_mux_153_nl;
  wire crc_mux_151_nl;
  wire crc_mux_149_nl;
  wire crc_mux_147_nl;
  wire crc_mux_145_nl;
  wire crc_mux_143_nl;
  wire crc_mux_141_nl;
  wire crc_mux_nl;
  wire crc_mux_167_nl;
  wire crc_mux_168_nl;
  wire crc_mux_169_nl;
  wire crc_mux_170_nl;
  wire crc_mux_171_nl;
  wire crc_mux_172_nl;
  wire crc_mux_173_nl;
  wire crc_mux_174_nl;
  wire crc_mux_175_nl;
  wire crc_mux_176_nl;
  wire crc_mux_177_nl;
  wire crc_mux_178_nl;
  wire crc_mux_179_nl;
  wire crc_mux_180_nl;
  wire crc_mux_181_nl;
  wire crc_mux_182_nl;
  wire crc_mux_183_nl;
  wire crc_mux_184_nl;
  wire crc_mux_185_nl;
  wire crc_mux_186_nl;
  wire crc_mux_187_nl;
  wire crc_mux_188_nl;
  wire crc_mux_189_nl;
  wire crc_mux_190_nl;
  wire crc_mux_191_nl;
  wire crc_mux_192_nl;
  wire crc_mux_193_nl;
  wire[8:0] for_acc_nl;
  wire[7:0] for_mux_2_nl;

  // Interconnect Declarations for Component Instantiations 
  wire [31:0] nl_crc32_core_out_rsci_inst_out_rsci_idat;
  assign nl_crc32_core_out_rsci_inst_out_rsci_idat = {out_rsci_idat_31 , out_rsci_idat_30
      , out_rsci_idat_29 , out_rsci_idat_28 , out_rsci_idat_27 , out_rsci_idat_26
      , out_rsci_idat_25 , out_rsci_idat_24 , out_rsci_idat_23 , out_rsci_idat_22
      , out_rsci_idat_21 , out_rsci_idat_20 , out_rsci_idat_19 , out_rsci_idat_18
      , out_rsci_idat_17 , out_rsci_idat_16 , out_rsci_idat_15 , out_rsci_idat_14
      , out_rsci_idat_13 , out_rsci_idat_12 , out_rsci_idat_11 , out_rsci_idat_10
      , out_rsci_idat_9 , out_rsci_idat_8 , out_rsci_idat_7 , out_rsci_idat_6 , out_rsci_idat_5
      , out_rsci_idat_4 , out_rsci_idat_3 , out_rsci_idat_2 , out_rsci_idat_1 , out_rsci_idat_0};
  crc32_core_in_rsci crc32_core_in_rsci_inst (
      .in_rsc_dat(in_rsc_dat),
      .in_rsc_vld(in_rsc_vld),
      .in_rsc_rdy(in_rsc_rdy),
      .in_rsci_oswt(reg_in_rsci_iswt0_cse),
      .in_rsci_wen_comp(in_rsci_wen_comp),
      .in_rsci_idat_mxwt(in_rsci_idat_mxwt)
    );
  crc32_core_out_rsci crc32_core_out_rsci_inst (
      .out_rsc_dat(out_rsc_dat),
      .out_rsc_vld(out_rsc_vld),
      .out_rsc_rdy(out_rsc_rdy),
      .out_rsci_oswt(reg_out_rsci_iswt0_cse),
      .out_rsci_wen_comp(out_rsci_wen_comp),
      .out_rsci_idat(nl_crc32_core_out_rsci_inst_out_rsci_idat[31:0])
    );
  crc32_core_staller crc32_core_staller_inst (
      .core_wen(core_wen),
      .in_rsci_wen_comp(in_rsci_wen_comp),
      .out_rsci_wen_comp(out_rsci_wen_comp)
    );
  crc32_core_core_fsm crc32_core_core_fsm_inst (
      .clk(clk),
      .rst(rst),
      .core_wen(core_wen),
      .fsm_output(fsm_output),
      .main_C_0_tr0(exit_for_sva_mx0),
      .for_C_0_tr0(exit_for_sva_mx0)
    );
  assign and_314_cse = core_wen & (~((fsm_output[0]) | (fsm_output[3]) | (~ exit_for_sva_mx0)));
  assign crc_mux_140_cse = MUX_s_1_2_2((~ crc_8_2_lpi_2_dfm_mx0), crc_8_2_lpi_2_dfm_mx0,
      not_tmp_4);
  assign for_acc_nl = $signed((z_out[7:0])) - $signed(size_val_sva);
  assign exit_for_sva_mx0 = MUX_s_1_2_2((~ (z_out[8])), (~ (readslicef_9_1_8(for_acc_nl))),
      fsm_output[2]);
  assign crc_5_4_lpi_2_dfm_mx0 = MUX_s_1_2_2((~ crc_8_1_sva), crc_8_1_sva, not_tmp_8);
  assign crc_8_2_lpi_2_dfm_mx0 = MUX_s_1_2_2((~ crc_9_1_sva), crc_9_1_sva, not_tmp_9);
  assign for_for_4_b_xor_tmp = (in_rsci_idat_mxwt[3]) ^ crc_3_1_sva;
  assign crc_8_3_lpi_2_dfm_mx0 = MUX_s_1_2_2((~ crc_9_2_lpi_2_dfm_mx0), crc_9_2_lpi_2_dfm_mx0,
      not_tmp_10);
  assign for_for_5_b_xor_tmp = (in_rsci_idat_mxwt[4]) ^ crc_4_1_sva;
  assign crc_8_4_lpi_2_dfm_mx0 = MUX_s_1_2_2((~ crc_9_3_lpi_2_dfm_mx0), crc_9_3_lpi_2_dfm_mx0,
      not_tmp_8);
  assign for_for_6_b_xor_tmp = (in_rsci_idat_mxwt[5]) ^ crc_5_1_sva;
  assign crc_8_5_lpi_2_dfm_mx0 = MUX_s_1_2_2((~ crc_9_4_lpi_2_dfm_mx0), crc_9_4_lpi_2_dfm_mx0,
      not_tmp_4);
  assign for_for_7_b_xor_tmp = (in_rsci_idat_mxwt[6]) ^ xor_cse_5;
  assign crc_8_6_lpi_2_dfm_mx0 = MUX_s_1_2_2((~ crc_9_5_lpi_2_dfm_mx0), crc_9_5_lpi_2_dfm_mx0,
      not_tmp_5);
  assign for_for_8_b_xor_tmp = (in_rsci_idat_mxwt[7]) ^ xor_cse_1;
  assign crc_9_6_lpi_2_dfm_mx0 = MUX_s_1_2_2((~ crc_14_1_sva), crc_14_1_sva, not_tmp_5);
  assign crc_9_7_lpi_2_dfm_mx0 = MUX_s_1_2_2((~ crc_15_1_sva), crc_15_1_sva, not_tmp_7);
  assign crc_9_lpi_2_dfm_mx0 = MUX_s_1_2_2((~ crc_15_2_lpi_2_dfm_mx0), crc_15_2_lpi_2_dfm_mx0,
      not_tmp_6);
  assign crc_15_3_lpi_2_dfm_mx0 = MUX_s_1_2_2((~ crc_17_1_sva), crc_17_1_sva, not_tmp_10);
  assign crc_15_4_lpi_2_dfm_mx0 = MUX_s_1_2_2((~ crc_18_1_sva), crc_18_1_sva, not_tmp_8);
  assign crc_15_5_lpi_2_dfm_mx0 = MUX_s_1_2_2((~ crc_19_1_sva), crc_19_1_sva, not_tmp_4);
  assign crc_19_2_lpi_2_dfm_mx0 = MUX_s_1_2_2((~ crc_20_1_sva), crc_20_1_sva, not_tmp_9);
  assign crc_19_3_lpi_2_dfm_mx0 = MUX_s_1_2_2((~ crc_20_2_lpi_2_dfm_mx0), crc_20_2_lpi_2_dfm_mx0,
      not_tmp_10);
  assign crc_19_4_lpi_2_dfm_mx0 = MUX_s_1_2_2((~ crc_20_3_lpi_2_dfm_mx0), crc_20_3_lpi_2_dfm_mx0,
      not_tmp_8);
  assign crc_19_5_lpi_2_dfm_mx0 = MUX_s_1_2_2((~ crc_20_4_lpi_2_dfm_mx0), crc_20_4_lpi_2_dfm_mx0,
      not_tmp_4);
  assign crc_20_5_lpi_2_dfm_mx0 = MUX_s_1_2_2((~ crc_21_4_lpi_2_dfm_mx0), crc_21_4_lpi_2_dfm_mx0,
      not_tmp_4);
  assign crc_20_6_lpi_2_dfm_mx0 = MUX_s_1_2_2((~ crc_21_5_lpi_2_dfm_mx0), crc_21_5_lpi_2_dfm_mx0,
      not_tmp_5);
  assign crc_20_7_lpi_2_dfm_mx0 = MUX_s_1_2_2((~ crc_21_6_lpi_2_dfm_mx0), crc_21_6_lpi_2_dfm_mx0,
      not_tmp_7);
  assign crc_20_lpi_2_dfm_mx0 = MUX_s_1_2_2((~ crc_21_7_lpi_2_dfm_mx0), crc_21_7_lpi_2_dfm_mx0,
      not_tmp_6);
  assign crc_21_lpi_2_dfm_mx0 = MUX_s_1_2_2((~ crc_23_6_lpi_2_dfm_mx0), crc_23_6_lpi_2_dfm_mx0,
      not_tmp_6);
  assign crc_23_7_lpi_2_dfm_mx0 = MUX_s_1_2_2((~ crc_24_6_lpi_2_dfm_mx0), crc_24_6_lpi_2_dfm_mx0,
      not_tmp_7);
  assign crc_24_7_lpi_2_dfm_mx0 = MUX_s_1_2_2((~ crc_26_5_lpi_2_dfm_mx0), crc_26_5_lpi_2_dfm_mx0,
      not_tmp_7);
  assign crc_24_lpi_2_dfm_mx0 = MUX_s_1_2_2((~ crc_26_6_lpi_2_dfm_mx0), crc_26_6_lpi_2_dfm_mx0,
      not_tmp_6);
  assign crc_26_7_lpi_2_dfm_mx0 = MUX_s_1_2_2((~ crc_27_6_lpi_2_dfm_mx0), crc_27_6_lpi_2_dfm_mx0,
      not_tmp_7);
  assign crc_27_7_lpi_2_dfm_mx0 = MUX_s_1_2_2((~ crc_29_5_lpi_2_dfm_mx0), crc_29_5_lpi_2_dfm_mx0,
      not_tmp_7);
  assign crc_27_lpi_2_dfm_mx0 = MUX_s_1_2_2((~ crc_29_6_lpi_2_dfm_mx0), crc_29_6_lpi_2_dfm_mx0,
      not_tmp_6);
  assign crc_29_7_lpi_2_dfm_mx0 = MUX_s_1_2_2((~ crc_30_6_lpi_2_dfm_mx0), crc_30_6_lpi_2_dfm_mx0,
      not_tmp_7);
  assign crc_30_7_lpi_2_dfm_mx0 = MUX_s_1_2_2((~ for_for_5_b_xor_tmp), for_for_5_b_xor_tmp,
      not_tmp_7);
  assign crc_30_lpi_2_dfm_mx0 = MUX_s_1_2_2((~ for_for_6_b_xor_tmp), for_for_6_b_xor_tmp,
      not_tmp_6);
  assign for_for_b_2_sva_1 = (in_rsci_idat_mxwt[1]) ^ crc_1_1_sva;
  assign crc_15_2_lpi_2_dfm_mx0 = MUX_s_1_2_2((~ crc_16_1_sva), crc_16_1_sva, not_tmp_9);
  assign crc_21_7_lpi_2_dfm_mx0 = MUX_s_1_2_2((~ crc_23_5_lpi_2_dfm_mx0), crc_23_5_lpi_2_dfm_mx0,
      not_tmp_7);
  assign crc_23_6_lpi_2_dfm_mx0 = MUX_s_1_2_2((~ crc_24_5_lpi_2_dfm_mx0), crc_24_5_lpi_2_dfm_mx0,
      not_tmp_5);
  assign crc_26_6_lpi_2_dfm_mx0 = MUX_s_1_2_2((~ crc_27_5_lpi_2_dfm_mx0), crc_27_5_lpi_2_dfm_mx0,
      not_tmp_5);
  assign crc_29_6_lpi_2_dfm_mx0 = MUX_s_1_2_2((~ crc_30_5_lpi_2_dfm_mx0), crc_30_5_lpi_2_dfm_mx0,
      not_tmp_5);
  assign for_for_b_1_sva_1 = (in_rsci_idat_mxwt[0]) ^ crc_0_1_sva;
  assign crc_21_6_lpi_2_dfm_mx0 = MUX_s_1_2_2((~ crc_23_4_lpi_2_dfm_mx0), crc_23_4_lpi_2_dfm_mx0,
      not_tmp_5);
  assign crc_23_5_lpi_2_dfm_mx0 = MUX_s_1_2_2((~ crc_24_4_lpi_2_dfm_mx0), crc_24_4_lpi_2_dfm_mx0,
      not_tmp_4);
  assign crc_24_6_lpi_2_dfm_mx0 = MUX_s_1_2_2((~ crc_26_4_lpi_2_dfm_mx0), crc_26_4_lpi_2_dfm_mx0,
      not_tmp_5);
  assign crc_26_5_lpi_2_dfm_mx0 = MUX_s_1_2_2((~ crc_27_4_lpi_2_dfm_mx0), crc_27_4_lpi_2_dfm_mx0,
      not_tmp_4);
  assign crc_27_6_lpi_2_dfm_mx0 = MUX_s_1_2_2((~ crc_29_4_lpi_2_dfm_mx0), crc_29_4_lpi_2_dfm_mx0,
      not_tmp_5);
  assign crc_29_5_lpi_2_dfm_mx0 = MUX_s_1_2_2((~ crc_30_4_lpi_2_dfm_mx0), crc_30_4_lpi_2_dfm_mx0,
      not_tmp_4);
  assign crc_30_6_lpi_2_dfm_mx0 = MUX_s_1_2_2((~ for_for_4_b_xor_tmp), for_for_4_b_xor_tmp,
      not_tmp_5);
  assign crc_9_5_lpi_2_dfm_mx0 = MUX_s_1_2_2((~ crc_13_1_sva), crc_13_1_sva, not_tmp_4);
  assign crc_21_5_lpi_2_dfm_mx0 = MUX_s_1_2_2((~ crc_23_3_lpi_2_dfm_mx0), crc_23_3_lpi_2_dfm_mx0,
      not_tmp_4);
  assign crc_23_4_lpi_2_dfm_mx0 = MUX_s_1_2_2((~ crc_24_3_lpi_2_dfm_mx0), crc_24_3_lpi_2_dfm_mx0,
      not_tmp_8);
  assign crc_24_5_lpi_2_dfm_mx0 = MUX_s_1_2_2((~ crc_26_3_lpi_2_dfm_mx0), crc_26_3_lpi_2_dfm_mx0,
      not_tmp_4);
  assign crc_26_4_lpi_2_dfm_mx0 = MUX_s_1_2_2((~ crc_27_3_lpi_2_dfm_mx0), crc_27_3_lpi_2_dfm_mx0,
      not_tmp_8);
  assign crc_27_5_lpi_2_dfm_mx0 = MUX_s_1_2_2((~ crc_29_3_lpi_2_dfm_mx0), crc_29_3_lpi_2_dfm_mx0,
      not_tmp_4);
  assign crc_29_4_lpi_2_dfm_mx0 = MUX_s_1_2_2((~ crc_30_3_lpi_2_dfm_mx0), crc_30_3_lpi_2_dfm_mx0,
      not_tmp_8);
  assign crc_30_5_lpi_2_dfm_mx0 = MUX_s_1_2_2((~ for_for_b_3_sva_1), for_for_b_3_sva_1,
      not_tmp_4);
  assign crc_9_4_lpi_2_dfm_mx0 = MUX_s_1_2_2((~ crc_12_1_sva), crc_12_1_sva, not_tmp_8);
  assign crc_20_4_lpi_2_dfm_mx0 = MUX_s_1_2_2((~ crc_21_3_lpi_2_dfm_mx0), crc_21_3_lpi_2_dfm_mx0,
      not_tmp_8);
  assign crc_21_4_lpi_2_dfm_mx0 = MUX_s_1_2_2((~ crc_23_2_lpi_2_dfm_mx0), crc_23_2_lpi_2_dfm_mx0,
      not_tmp_8);
  assign crc_23_3_lpi_2_dfm_mx0 = MUX_s_1_2_2((~ crc_24_2_lpi_2_dfm_mx0), crc_24_2_lpi_2_dfm_mx0,
      not_tmp_10);
  assign crc_24_4_lpi_2_dfm_mx0 = MUX_s_1_2_2((~ crc_26_2_lpi_2_dfm_mx0), crc_26_2_lpi_2_dfm_mx0,
      not_tmp_8);
  assign crc_26_3_lpi_2_dfm_mx0 = MUX_s_1_2_2((~ crc_27_2_lpi_2_dfm_mx0), crc_27_2_lpi_2_dfm_mx0,
      not_tmp_10);
  assign crc_27_4_lpi_2_dfm_mx0 = MUX_s_1_2_2((~ crc_29_2_lpi_2_dfm_mx0), crc_29_2_lpi_2_dfm_mx0,
      not_tmp_8);
  assign crc_29_3_lpi_2_dfm_mx0 = MUX_s_1_2_2((~ crc_30_2_lpi_2_dfm_mx0), crc_30_2_lpi_2_dfm_mx0,
      not_tmp_10);
  assign crc_30_4_lpi_2_dfm_mx0 = MUX_s_1_2_2((~ for_for_b_2_sva_1), for_for_b_2_sva_1,
      not_tmp_8);
  assign for_for_b_3_sva_1 = (in_rsci_idat_mxwt[2]) ^ crc_2_1_sva;
  assign crc_9_3_lpi_2_dfm_mx0 = MUX_s_1_2_2((~ crc_11_1_sva), crc_11_1_sva, not_tmp_10);
  assign crc_20_3_lpi_2_dfm_mx0 = MUX_s_1_2_2((~ crc_21_2_lpi_2_dfm_mx0), crc_21_2_lpi_2_dfm_mx0,
      not_tmp_10);
  assign crc_21_3_lpi_2_dfm_mx0 = MUX_s_1_2_2((~ crc_23_1_sva), crc_23_1_sva, not_tmp_10);
  assign crc_23_2_lpi_2_dfm_mx0 = MUX_s_1_2_2((~ crc_24_1_sva), crc_24_1_sva, not_tmp_9);
  assign crc_24_3_lpi_2_dfm_mx0 = MUX_s_1_2_2((~ crc_26_1_sva), crc_26_1_sva, not_tmp_10);
  assign crc_26_2_lpi_2_dfm_mx0 = MUX_s_1_2_2((~ crc_27_1_sva), crc_27_1_sva, not_tmp_9);
  assign crc_27_3_lpi_2_dfm_mx0 = MUX_s_1_2_2((~ crc_29_1_sva), crc_29_1_sva, not_tmp_10);
  assign crc_29_2_lpi_2_dfm_mx0 = MUX_s_1_2_2((~ crc_30_1_sva), crc_30_1_sva, not_tmp_9);
  assign crc_30_3_lpi_2_dfm_mx0 = MUX_s_1_2_2((~ for_for_b_1_sva_1), for_for_b_1_sva_1,
      not_tmp_10);
  assign crc_9_2_lpi_2_dfm_mx0 = MUX_s_1_2_2((~ crc_10_1_sva), crc_10_1_sva, not_tmp_9);
  assign crc_20_2_lpi_2_dfm_mx0 = MUX_s_1_2_2((~ crc_21_1_sva), crc_21_1_sva, not_tmp_9);
  assign crc_21_2_lpi_2_dfm_mx0 = MUX_s_1_2_2((~ crc_22_1_sva), crc_22_1_sva, not_tmp_9);
  assign crc_24_2_lpi_2_dfm_mx0 = MUX_s_1_2_2((~ crc_25_1_sva), crc_25_1_sva, not_tmp_9);
  assign crc_27_2_lpi_2_dfm_mx0 = MUX_s_1_2_2((~ crc_28_1_sva), crc_28_1_sva, not_tmp_9);
  assign crc_30_2_lpi_2_dfm_mx0 = MUX_s_1_2_2((~ crc_31_1_sva), crc_31_1_sva, not_tmp_9);
  assign or_tmp_32 = exit_for_sva_mx0 & ((fsm_output[2:1]!=2'b00));
  assign or_tmp_40 = not_tmp_3 & (fsm_output[2]);
  assign or_tmp_52 = not_tmp_5 & (fsm_output[2]);
  assign or_tmp_56 = not_tmp_6 & (fsm_output[2]);
  assign or_tmp_60 = not_tmp_7 & (fsm_output[2]);
  assign xor_cse_1 = MUX_s_1_2_2(crc_7_1_sva, (~ crc_7_1_sva), for_for_b_2_sva_1);
  assign not_tmp_3 = ~((in_rsci_idat_mxwt[7]) ^ xor_cse_1);
  assign not_tmp_4 = ~((in_rsci_idat_mxwt[3]) ^ crc_3_1_sva);
  assign not_tmp_5 = ~((in_rsci_idat_mxwt[4]) ^ crc_4_1_sva);
  assign xor_cse_5 = MUX_s_1_2_2(crc_6_1_sva, (~ crc_6_1_sva), for_for_b_1_sva_1);
  assign not_tmp_6 = ~((in_rsci_idat_mxwt[6]) ^ xor_cse_5);
  assign not_tmp_7 = ~((in_rsci_idat_mxwt[5]) ^ crc_5_1_sva);
  assign not_tmp_8 = ~((in_rsci_idat_mxwt[2]) ^ crc_2_1_sva);
  assign not_tmp_9 = ~((in_rsci_idat_mxwt[0]) ^ crc_0_1_sva);
  assign not_tmp_10 = ~((in_rsci_idat_mxwt[1]) ^ crc_1_1_sva);
  always @(posedge clk) begin
    if ( rst ) begin
      out_rsci_idat_0 <= 1'b0;
      out_rsci_idat_1 <= 1'b0;
      out_rsci_idat_2 <= 1'b0;
      out_rsci_idat_3 <= 1'b0;
      out_rsci_idat_4 <= 1'b0;
      out_rsci_idat_5 <= 1'b0;
      out_rsci_idat_6 <= 1'b0;
      out_rsci_idat_7 <= 1'b0;
      out_rsci_idat_8 <= 1'b0;
      out_rsci_idat_9 <= 1'b0;
      out_rsci_idat_10 <= 1'b0;
      out_rsci_idat_11 <= 1'b0;
      out_rsci_idat_12 <= 1'b0;
      out_rsci_idat_13 <= 1'b0;
      out_rsci_idat_14 <= 1'b0;
      out_rsci_idat_15 <= 1'b0;
      out_rsci_idat_16 <= 1'b0;
      out_rsci_idat_17 <= 1'b0;
      out_rsci_idat_18 <= 1'b0;
      out_rsci_idat_19 <= 1'b0;
      out_rsci_idat_20 <= 1'b0;
      out_rsci_idat_21 <= 1'b0;
      out_rsci_idat_22 <= 1'b0;
      out_rsci_idat_23 <= 1'b0;
      out_rsci_idat_24 <= 1'b0;
      out_rsci_idat_25 <= 1'b0;
      out_rsci_idat_26 <= 1'b0;
      out_rsci_idat_27 <= 1'b0;
      out_rsci_idat_28 <= 1'b0;
      out_rsci_idat_29 <= 1'b0;
      out_rsci_idat_30 <= 1'b0;
      out_rsci_idat_31 <= 1'b0;
    end
    else if ( and_314_cse ) begin
      out_rsci_idat_0 <= ~(crc_5_4_lpi_2_dfm_mx0 | (~ (fsm_output[2])));
      out_rsci_idat_1 <= ~(crc_mux_140_cse | (~ (fsm_output[2])));
      out_rsci_idat_2 <= ~(crc_mux_142_nl | (~ (fsm_output[2])));
      out_rsci_idat_3 <= ~(crc_mux_144_nl | (~ (fsm_output[2])));
      out_rsci_idat_4 <= ~(crc_mux_146_nl | (~ (fsm_output[2])));
      out_rsci_idat_5 <= ~(crc_mux_148_nl | (~ (fsm_output[2])));
      out_rsci_idat_6 <= ~(crc_mux_150_nl | (~ (fsm_output[2])));
      out_rsci_idat_7 <= ~(crc_mux_152_nl | (~ (fsm_output[2])));
      out_rsci_idat_8 <= ~(crc_mux_154_nl | (~ (fsm_output[2])));
      out_rsci_idat_9 <= ~(crc_mux_156_nl | (~ (fsm_output[2])));
      out_rsci_idat_10 <= ~(crc_15_4_lpi_2_dfm_mx0 | (~ (fsm_output[2])));
      out_rsci_idat_11 <= ~(crc_15_5_lpi_2_dfm_mx0 | (~ (fsm_output[2])));
      out_rsci_idat_12 <= ~(crc_mux_160_nl | (~ (fsm_output[2])));
      out_rsci_idat_13 <= ~(crc_mux_162_nl | (~ (fsm_output[2])));
      out_rsci_idat_14 <= ~(crc_mux_164_nl | (~ (fsm_output[2])));
      out_rsci_idat_15 <= ~(crc_mux_166_nl | (~ (fsm_output[2])));
      out_rsci_idat_16 <= ~(crc_mux_165_nl | (~ (fsm_output[2])));
      out_rsci_idat_17 <= ~(crc_mux_163_nl | (~ (fsm_output[2])));
      out_rsci_idat_18 <= ~(crc_mux_161_nl | (~ (fsm_output[2])));
      out_rsci_idat_19 <= ~(crc_mux_159_nl | (~ (fsm_output[2])));
      out_rsci_idat_20 <= ~(crc_mux_158_nl | (~ (fsm_output[2])));
      out_rsci_idat_21 <= ~(crc_mux_157_nl | (~ (fsm_output[2])));
      out_rsci_idat_22 <= ~(crc_mux_155_nl | (~ (fsm_output[2])));
      out_rsci_idat_23 <= ~(crc_mux_153_nl | (~ (fsm_output[2])));
      out_rsci_idat_24 <= ~(crc_mux_151_nl | (~ (fsm_output[2])));
      out_rsci_idat_25 <= ~(crc_mux_149_nl | (~ (fsm_output[2])));
      out_rsci_idat_26 <= ~(crc_mux_147_nl | (~ (fsm_output[2])));
      out_rsci_idat_27 <= ~(crc_mux_145_nl | (~ (fsm_output[2])));
      out_rsci_idat_28 <= ~(crc_mux_143_nl | (~ (fsm_output[2])));
      out_rsci_idat_29 <= ~(crc_mux_141_nl | (~ (fsm_output[2])));
      out_rsci_idat_30 <= ~(crc_mux_nl | (~ (fsm_output[2])));
      out_rsci_idat_31 <= ~(for_for_8_b_xor_tmp | (~ (fsm_output[2])));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_out_rsci_iswt0_cse <= 1'b0;
      reg_in_rsci_iswt0_cse <= 1'b0;
      crc_31_1_sva <= 1'b0;
      crc_0_1_sva <= 1'b0;
      crc_30_1_sva <= 1'b0;
      crc_1_1_sva <= 1'b0;
      crc_29_1_sva <= 1'b0;
      crc_2_1_sva <= 1'b0;
      crc_28_1_sva <= 1'b0;
      crc_3_1_sva <= 1'b0;
      crc_27_1_sva <= 1'b0;
      crc_4_1_sva <= 1'b0;
      crc_26_1_sva <= 1'b0;
      crc_5_1_sva <= 1'b0;
      crc_25_1_sva <= 1'b0;
      crc_6_1_sva <= 1'b0;
      crc_24_1_sva <= 1'b0;
      crc_7_1_sva <= 1'b0;
      crc_23_1_sva <= 1'b0;
      crc_8_1_sva <= 1'b0;
      crc_22_1_sva <= 1'b0;
      crc_9_1_sva <= 1'b0;
      crc_21_1_sva <= 1'b0;
      crc_10_1_sva <= 1'b0;
      crc_20_1_sva <= 1'b0;
      crc_11_1_sva <= 1'b0;
      crc_19_1_sva <= 1'b0;
      crc_12_1_sva <= 1'b0;
      crc_18_1_sva <= 1'b0;
      crc_13_1_sva <= 1'b0;
      crc_17_1_sva <= 1'b0;
      crc_14_1_sva <= 1'b0;
      crc_16_1_sva <= 1'b0;
      crc_15_1_sva <= 1'b0;
      for_i_sva <= 8'b00000000;
    end
    else if ( core_wen ) begin
      reg_out_rsci_iswt0_cse <= or_tmp_32;
      reg_in_rsci_iswt0_cse <= ~ or_tmp_32;
      crc_31_1_sva <= for_for_8_b_xor_tmp | (~ (fsm_output[2]));
      crc_0_1_sva <= crc_5_4_lpi_2_dfm_mx0 | (~ (fsm_output[2]));
      crc_30_1_sva <= crc_mux_167_nl | (~ (fsm_output[2]));
      crc_1_1_sva <= crc_mux_140_cse | (~ (fsm_output[2]));
      crc_29_1_sva <= crc_mux_168_nl | (~ (fsm_output[2]));
      crc_2_1_sva <= crc_mux_169_nl | (~ (fsm_output[2]));
      crc_28_1_sva <= crc_mux_170_nl | (~ (fsm_output[2]));
      crc_3_1_sva <= crc_mux_171_nl | (~ (fsm_output[2]));
      crc_27_1_sva <= crc_mux_172_nl | (~ (fsm_output[2]));
      crc_4_1_sva <= crc_mux_173_nl | (~ (fsm_output[2]));
      crc_26_1_sva <= crc_mux_174_nl | (~ (fsm_output[2]));
      crc_5_1_sva <= crc_mux_175_nl | (~ (fsm_output[2]));
      crc_25_1_sva <= crc_mux_176_nl | (~ (fsm_output[2]));
      crc_6_1_sva <= crc_mux_177_nl | (~ (fsm_output[2]));
      crc_24_1_sva <= crc_mux_178_nl | (~ (fsm_output[2]));
      crc_7_1_sva <= crc_mux_179_nl | (~ (fsm_output[2]));
      crc_23_1_sva <= crc_mux_180_nl | (~ (fsm_output[2]));
      crc_8_1_sva <= crc_mux_181_nl | (~ (fsm_output[2]));
      crc_22_1_sva <= crc_mux_182_nl | (~ (fsm_output[2]));
      crc_9_1_sva <= crc_mux_183_nl | (~ (fsm_output[2]));
      crc_21_1_sva <= crc_mux_184_nl | (~ (fsm_output[2]));
      crc_10_1_sva <= crc_15_4_lpi_2_dfm_mx0 | (~ (fsm_output[2]));
      crc_20_1_sva <= crc_mux_185_nl | (~ (fsm_output[2]));
      crc_11_1_sva <= crc_15_5_lpi_2_dfm_mx0 | (~ (fsm_output[2]));
      crc_19_1_sva <= crc_mux_186_nl | (~ (fsm_output[2]));
      crc_12_1_sva <= crc_mux_187_nl | (~ (fsm_output[2]));
      crc_18_1_sva <= crc_mux_188_nl | (~ (fsm_output[2]));
      crc_13_1_sva <= crc_mux_189_nl | (~ (fsm_output[2]));
      crc_17_1_sva <= crc_mux_190_nl | (~ (fsm_output[2]));
      crc_14_1_sva <= crc_mux_191_nl | (~ (fsm_output[2]));
      crc_16_1_sva <= crc_mux_192_nl | (~ (fsm_output[2]));
      crc_15_1_sva <= crc_mux_193_nl | (~ (fsm_output[2]));
      for_i_sva <= MUX_v_8_2_2(8'b00000000, (z_out[7:0]), (fsm_output[2]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      size_val_sva <= 8'b00000000;
    end
    else if ( core_wen & (~ (fsm_output[2])) ) begin
      size_val_sva <= in_rsci_idat_mxwt;
    end
  end
  assign crc_mux_142_nl = MUX_s_1_2_2((~ crc_8_3_lpi_2_dfm_mx0), crc_8_3_lpi_2_dfm_mx0,
      or_tmp_52);
  assign crc_mux_144_nl = MUX_s_1_2_2((~ crc_8_4_lpi_2_dfm_mx0), crc_8_4_lpi_2_dfm_mx0,
      or_tmp_60);
  assign crc_mux_146_nl = MUX_s_1_2_2((~ crc_8_5_lpi_2_dfm_mx0), crc_8_5_lpi_2_dfm_mx0,
      or_tmp_56);
  assign crc_mux_148_nl = MUX_s_1_2_2((~ crc_8_6_lpi_2_dfm_mx0), crc_8_6_lpi_2_dfm_mx0,
      or_tmp_40);
  assign crc_mux_150_nl = MUX_s_1_2_2((~ crc_9_6_lpi_2_dfm_mx0), crc_9_6_lpi_2_dfm_mx0,
      or_tmp_60);
  assign crc_mux_152_nl = MUX_s_1_2_2((~ crc_9_7_lpi_2_dfm_mx0), crc_9_7_lpi_2_dfm_mx0,
      or_tmp_56);
  assign crc_mux_154_nl = MUX_s_1_2_2((~ crc_9_lpi_2_dfm_mx0), crc_9_lpi_2_dfm_mx0,
      or_tmp_40);
  assign crc_mux_156_nl = MUX_s_1_2_2((~ crc_15_3_lpi_2_dfm_mx0), crc_15_3_lpi_2_dfm_mx0,
      or_tmp_40);
  assign crc_mux_160_nl = MUX_s_1_2_2((~ crc_19_2_lpi_2_dfm_mx0), crc_19_2_lpi_2_dfm_mx0,
      or_tmp_52);
  assign crc_mux_162_nl = MUX_s_1_2_2((~ crc_19_3_lpi_2_dfm_mx0), crc_19_3_lpi_2_dfm_mx0,
      or_tmp_60);
  assign crc_mux_164_nl = MUX_s_1_2_2((~ crc_19_4_lpi_2_dfm_mx0), crc_19_4_lpi_2_dfm_mx0,
      or_tmp_56);
  assign crc_mux_166_nl = MUX_s_1_2_2((~ crc_19_5_lpi_2_dfm_mx0), crc_19_5_lpi_2_dfm_mx0,
      or_tmp_40);
  assign crc_mux_165_nl = MUX_s_1_2_2((~ crc_20_5_lpi_2_dfm_mx0), crc_20_5_lpi_2_dfm_mx0,
      or_tmp_52);
  assign crc_mux_163_nl = MUX_s_1_2_2((~ crc_20_6_lpi_2_dfm_mx0), crc_20_6_lpi_2_dfm_mx0,
      or_tmp_60);
  assign crc_mux_161_nl = MUX_s_1_2_2((~ crc_20_7_lpi_2_dfm_mx0), crc_20_7_lpi_2_dfm_mx0,
      or_tmp_56);
  assign crc_mux_159_nl = MUX_s_1_2_2((~ crc_20_lpi_2_dfm_mx0), crc_20_lpi_2_dfm_mx0,
      or_tmp_40);
  assign crc_mux_158_nl = MUX_s_1_2_2((~ crc_21_lpi_2_dfm_mx0), crc_21_lpi_2_dfm_mx0,
      or_tmp_40);
  assign crc_mux_157_nl = MUX_s_1_2_2((~ crc_23_7_lpi_2_dfm_mx0), crc_23_7_lpi_2_dfm_mx0,
      or_tmp_40);
  assign crc_mux_155_nl = MUX_s_1_2_2((~ crc_24_7_lpi_2_dfm_mx0), crc_24_7_lpi_2_dfm_mx0,
      or_tmp_56);
  assign crc_mux_153_nl = MUX_s_1_2_2((~ crc_24_lpi_2_dfm_mx0), crc_24_lpi_2_dfm_mx0,
      or_tmp_40);
  assign crc_mux_151_nl = MUX_s_1_2_2((~ crc_26_7_lpi_2_dfm_mx0), crc_26_7_lpi_2_dfm_mx0,
      or_tmp_40);
  assign crc_mux_149_nl = MUX_s_1_2_2((~ crc_27_7_lpi_2_dfm_mx0), crc_27_7_lpi_2_dfm_mx0,
      or_tmp_56);
  assign crc_mux_147_nl = MUX_s_1_2_2((~ crc_27_lpi_2_dfm_mx0), crc_27_lpi_2_dfm_mx0,
      or_tmp_40);
  assign crc_mux_145_nl = MUX_s_1_2_2((~ crc_29_7_lpi_2_dfm_mx0), crc_29_7_lpi_2_dfm_mx0,
      or_tmp_40);
  assign crc_mux_143_nl = MUX_s_1_2_2((~ crc_30_7_lpi_2_dfm_mx0), crc_30_7_lpi_2_dfm_mx0,
      or_tmp_56);
  assign crc_mux_141_nl = MUX_s_1_2_2((~ crc_30_lpi_2_dfm_mx0), crc_30_lpi_2_dfm_mx0,
      or_tmp_40);
  assign crc_mux_nl = MUX_s_1_2_2((~ for_for_7_b_xor_tmp), for_for_7_b_xor_tmp, or_tmp_40);
  assign crc_mux_167_nl = MUX_s_1_2_2((~ for_for_7_b_xor_tmp), for_for_7_b_xor_tmp,
      not_tmp_3);
  assign crc_mux_168_nl = MUX_s_1_2_2((~ crc_30_lpi_2_dfm_mx0), crc_30_lpi_2_dfm_mx0,
      not_tmp_3);
  assign crc_mux_169_nl = MUX_s_1_2_2((~ crc_8_3_lpi_2_dfm_mx0), crc_8_3_lpi_2_dfm_mx0,
      not_tmp_5);
  assign crc_mux_170_nl = MUX_s_1_2_2((~ crc_30_7_lpi_2_dfm_mx0), crc_30_7_lpi_2_dfm_mx0,
      not_tmp_6);
  assign crc_mux_171_nl = MUX_s_1_2_2((~ crc_8_4_lpi_2_dfm_mx0), crc_8_4_lpi_2_dfm_mx0,
      not_tmp_7);
  assign crc_mux_172_nl = MUX_s_1_2_2((~ crc_29_7_lpi_2_dfm_mx0), crc_29_7_lpi_2_dfm_mx0,
      not_tmp_3);
  assign crc_mux_173_nl = MUX_s_1_2_2((~ crc_8_5_lpi_2_dfm_mx0), crc_8_5_lpi_2_dfm_mx0,
      not_tmp_6);
  assign crc_mux_174_nl = MUX_s_1_2_2((~ crc_27_lpi_2_dfm_mx0), crc_27_lpi_2_dfm_mx0,
      not_tmp_3);
  assign crc_mux_175_nl = MUX_s_1_2_2((~ crc_8_6_lpi_2_dfm_mx0), crc_8_6_lpi_2_dfm_mx0,
      not_tmp_3);
  assign crc_mux_176_nl = MUX_s_1_2_2((~ crc_27_7_lpi_2_dfm_mx0), crc_27_7_lpi_2_dfm_mx0,
      not_tmp_6);
  assign crc_mux_177_nl = MUX_s_1_2_2((~ crc_9_6_lpi_2_dfm_mx0), crc_9_6_lpi_2_dfm_mx0,
      not_tmp_7);
  assign crc_mux_178_nl = MUX_s_1_2_2((~ crc_26_7_lpi_2_dfm_mx0), crc_26_7_lpi_2_dfm_mx0,
      not_tmp_3);
  assign crc_mux_179_nl = MUX_s_1_2_2((~ crc_9_7_lpi_2_dfm_mx0), crc_9_7_lpi_2_dfm_mx0,
      not_tmp_6);
  assign crc_mux_180_nl = MUX_s_1_2_2((~ crc_24_lpi_2_dfm_mx0), crc_24_lpi_2_dfm_mx0,
      not_tmp_3);
  assign crc_mux_181_nl = MUX_s_1_2_2((~ crc_9_lpi_2_dfm_mx0), crc_9_lpi_2_dfm_mx0,
      not_tmp_3);
  assign crc_mux_182_nl = MUX_s_1_2_2((~ crc_24_7_lpi_2_dfm_mx0), crc_24_7_lpi_2_dfm_mx0,
      not_tmp_6);
  assign crc_mux_183_nl = MUX_s_1_2_2((~ crc_15_3_lpi_2_dfm_mx0), crc_15_3_lpi_2_dfm_mx0,
      not_tmp_3);
  assign crc_mux_184_nl = MUX_s_1_2_2((~ crc_23_7_lpi_2_dfm_mx0), crc_23_7_lpi_2_dfm_mx0,
      not_tmp_3);
  assign crc_mux_185_nl = MUX_s_1_2_2((~ crc_21_lpi_2_dfm_mx0), crc_21_lpi_2_dfm_mx0,
      not_tmp_3);
  assign crc_mux_186_nl = MUX_s_1_2_2((~ crc_20_lpi_2_dfm_mx0), crc_20_lpi_2_dfm_mx0,
      not_tmp_3);
  assign crc_mux_187_nl = MUX_s_1_2_2((~ crc_19_2_lpi_2_dfm_mx0), crc_19_2_lpi_2_dfm_mx0,
      not_tmp_5);
  assign crc_mux_188_nl = MUX_s_1_2_2((~ crc_20_7_lpi_2_dfm_mx0), crc_20_7_lpi_2_dfm_mx0,
      not_tmp_6);
  assign crc_mux_189_nl = MUX_s_1_2_2((~ crc_19_3_lpi_2_dfm_mx0), crc_19_3_lpi_2_dfm_mx0,
      not_tmp_7);
  assign crc_mux_190_nl = MUX_s_1_2_2((~ crc_20_6_lpi_2_dfm_mx0), crc_20_6_lpi_2_dfm_mx0,
      not_tmp_7);
  assign crc_mux_191_nl = MUX_s_1_2_2((~ crc_19_4_lpi_2_dfm_mx0), crc_19_4_lpi_2_dfm_mx0,
      not_tmp_6);
  assign crc_mux_192_nl = MUX_s_1_2_2((~ crc_20_5_lpi_2_dfm_mx0), crc_20_5_lpi_2_dfm_mx0,
      not_tmp_5);
  assign crc_mux_193_nl = MUX_s_1_2_2((~ crc_19_5_lpi_2_dfm_mx0), crc_19_5_lpi_2_dfm_mx0,
      not_tmp_3);
  assign for_mux_2_nl = MUX_v_8_2_2((~ in_rsci_idat_mxwt), for_i_sva, fsm_output[2]);
  assign nl_z_out = conv_s2u_8_9(for_mux_2_nl) + 9'b000000001;
  assign z_out = nl_z_out[8:0];

  function automatic  MUX_s_1_2_2;
    input  input_0;
    input  input_1;
    input  sel;
    reg  result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [7:0] MUX_v_8_2_2;
    input [7:0] input_0;
    input [7:0] input_1;
    input  sel;
    reg [7:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_8_2_2 = result;
  end
  endfunction


  function automatic [0:0] readslicef_9_1_8;
    input [8:0] vector;
    reg [8:0] tmp;
  begin
    tmp = vector >> 8;
    readslicef_9_1_8 = tmp[0:0];
  end
  endfunction


  function automatic [8:0] conv_s2u_8_9 ;
    input [7:0]  vector ;
  begin
    conv_s2u_8_9 = {vector[7], vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    crc32
// ------------------------------------------------------------------


module crc32 (
  clk, rst, in_rsc_dat, in_rsc_vld, in_rsc_rdy, out_rsc_dat, out_rsc_vld, out_rsc_rdy
);
  input clk;
  input rst;
  input [7:0] in_rsc_dat;
  input in_rsc_vld;
  output in_rsc_rdy;
  output [31:0] out_rsc_dat;
  output out_rsc_vld;
  input out_rsc_rdy;



  // Interconnect Declarations for Component Instantiations 
  crc32_core crc32_core_inst (
      .clk(clk),
      .rst(rst),
      .in_rsc_dat(in_rsc_dat),
      .in_rsc_vld(in_rsc_vld),
      .in_rsc_rdy(in_rsc_rdy),
      .out_rsc_dat(out_rsc_dat),
      .out_rsc_vld(out_rsc_vld),
      .out_rsc_rdy(out_rsc_rdy)
    );
endmodule




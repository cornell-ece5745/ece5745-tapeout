magic
tech sky130A
magscale 1 2
timestamp 1655493482
<< obsli1 >>
rect 1104 2159 138828 137649
<< obsm1 >>
rect 1104 2128 138828 137680
<< metal2 >>
rect 14002 139200 14058 140000
rect 41970 139200 42026 140000
rect 69938 139200 69994 140000
rect 97998 139200 98054 140000
rect 125966 139200 126022 140000
rect 9954 0 10010 800
rect 29918 0 29974 800
rect 49882 0 49938 800
rect 69938 0 69994 800
rect 89902 0 89958 800
rect 109958 0 110014 800
rect 129922 0 129978 800
<< obsm2 >>
rect 1398 139144 13946 139346
rect 14114 139144 41914 139346
rect 42082 139144 69882 139346
rect 70050 139144 97942 139346
rect 98110 139144 125910 139346
rect 126078 139144 138166 139346
rect 1398 856 138166 139144
rect 1398 800 9898 856
rect 10066 800 29862 856
rect 30030 800 49826 856
rect 49994 800 69882 856
rect 70050 800 89846 856
rect 90014 800 109902 856
rect 110070 800 129866 856
rect 130034 800 138166 856
<< metal3 >>
rect 0 122272 800 122392
rect 139200 104864 140000 104984
rect 0 87320 800 87440
rect 0 52368 800 52488
rect 139200 34960 140000 35080
rect 0 17416 800 17536
<< obsm3 >>
rect 800 122472 139200 137665
rect 880 122192 139200 122472
rect 800 105064 139200 122192
rect 800 104784 139120 105064
rect 800 87520 139200 104784
rect 880 87240 139200 87520
rect 800 52568 139200 87240
rect 880 52288 139200 52568
rect 800 35160 139200 52288
rect 800 34880 139120 35160
rect 800 17616 139200 34880
rect 880 17336 139200 17616
rect 800 2143 139200 17336
<< metal4 >>
rect 4208 2128 4528 137680
rect 19568 2128 19888 137680
rect 34928 2128 35248 137680
rect 50288 2128 50608 137680
rect 65648 2128 65968 137680
rect 81008 2128 81328 137680
rect 96368 2128 96688 137680
rect 111728 2128 112048 137680
rect 127088 2128 127408 137680
<< obsm4 >>
rect 61515 33627 61581 61029
<< labels >>
rlabel metal2 s 49882 0 49938 800 6 adapter_parity
port 1 nsew signal output
rlabel metal2 s 69938 0 69994 800 6 ap_en
port 2 nsew signal output
rlabel metal2 s 14002 139200 14058 140000 6 clk
port 3 nsew signal input
rlabel metal2 s 41970 139200 42026 140000 6 clk_en
port 4 nsew signal output
rlabel metal3 s 0 87320 800 87440 6 cs_en
port 5 nsew signal output
rlabel metal2 s 9954 0 10010 800 6 loopthrough_sel
port 6 nsew signal input
rlabel metal2 s 89902 0 89958 800 6 lt_sel_en
port 7 nsew signal output
rlabel metal2 s 29918 0 29974 800 6 minion_parity
port 8 nsew signal output
rlabel metal2 s 109958 0 110014 800 6 miso_en
port 9 nsew signal output
rlabel metal2 s 125966 139200 126022 140000 6 mosi_en
port 10 nsew signal output
rlabel metal2 s 129922 0 129978 800 6 mp_en
port 11 nsew signal output
rlabel metal2 s 69938 139200 69994 140000 6 reset
port 12 nsew signal input
rlabel metal2 s 97998 139200 98054 140000 6 reset_en
port 13 nsew signal output
rlabel metal3 s 0 122272 800 122392 6 sclk_en
port 14 nsew signal output
rlabel metal3 s 139200 34960 140000 35080 6 spi_min_cs
port 15 nsew signal input
rlabel metal3 s 0 52368 800 52488 6 spi_min_miso
port 16 nsew signal output
rlabel metal3 s 0 17416 800 17536 6 spi_min_mosi
port 17 nsew signal input
rlabel metal3 s 139200 104864 140000 104984 6 spi_min_sclk
port 18 nsew signal input
rlabel metal4 s 4208 2128 4528 137680 6 vccd1
port 19 nsew power input
rlabel metal4 s 34928 2128 35248 137680 6 vccd1
port 19 nsew power input
rlabel metal4 s 65648 2128 65968 137680 6 vccd1
port 19 nsew power input
rlabel metal4 s 96368 2128 96688 137680 6 vccd1
port 19 nsew power input
rlabel metal4 s 127088 2128 127408 137680 6 vccd1
port 19 nsew power input
rlabel metal4 s 19568 2128 19888 137680 6 vssd1
port 20 nsew ground input
rlabel metal4 s 50288 2128 50608 137680 6 vssd1
port 20 nsew ground input
rlabel metal4 s 81008 2128 81328 137680 6 vssd1
port 20 nsew ground input
rlabel metal4 s 111728 2128 112048 137680 6 vssd1
port 20 nsew ground input
<< properties >>
string FIXED_BBOX 0 0 140000 140000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 12680174
string GDS_FILE /home/acm289/ece5745-tapeout/openlane/project-group15/runs/project-group15/results/finishing/grp_15_SPI_TapeOutBlockRTL_32bits_5entries.magic.gds
string GDS_START 642594
<< end >>


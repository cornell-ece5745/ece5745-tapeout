magic
tech sky130A
magscale 1 2
timestamp 1655493474
<< obsli1 >>
rect 1104 2159 138828 137649
<< obsm1 >>
rect 1104 2128 138828 137680
<< metal2 >>
rect 11610 139200 11666 140000
rect 34886 139200 34942 140000
rect 58254 139200 58310 140000
rect 81622 139200 81678 140000
rect 104898 139200 104954 140000
rect 128266 139200 128322 140000
rect 11610 0 11666 800
rect 34886 0 34942 800
rect 58254 0 58310 800
rect 81622 0 81678 800
rect 104898 0 104954 800
rect 128266 0 128322 800
<< obsm2 >>
rect 1398 139144 11554 139346
rect 11722 139144 34830 139346
rect 34998 139144 58198 139346
rect 58366 139144 81566 139346
rect 81734 139144 104842 139346
rect 105010 139144 128210 139346
rect 128378 139144 138166 139346
rect 1398 856 138166 139144
rect 1398 800 11554 856
rect 11722 800 34830 856
rect 34998 800 58198 856
rect 58366 800 81566 856
rect 81734 800 104842 856
rect 105010 800 128210 856
rect 128378 800 138166 856
<< metal3 >>
rect 0 116560 800 116680
rect 139200 116560 140000 116680
rect 0 69912 800 70032
rect 139200 69912 140000 70032
rect 0 23264 800 23384
rect 139200 23264 140000 23384
<< obsm3 >>
rect 800 116760 139200 137665
rect 880 116480 139120 116760
rect 800 70112 139200 116480
rect 880 69832 139120 70112
rect 800 23464 139200 69832
rect 880 23184 139120 23464
rect 800 2143 139200 23184
<< metal4 >>
rect 4208 2128 4528 137680
rect 19568 2128 19888 137680
rect 34928 2128 35248 137680
rect 50288 2128 50608 137680
rect 65648 2128 65968 137680
rect 81008 2128 81328 137680
rect 96368 2128 96688 137680
rect 111728 2128 112048 137680
rect 127088 2128 127408 137680
<< obsm4 >>
rect 77891 23699 80928 117333
rect 81408 23699 90837 117333
<< labels >>
rlabel metal3 s 139200 116560 140000 116680 6 adapter_parity
port 1 nsew signal output
rlabel metal3 s 0 23264 800 23384 6 ap_en
port 2 nsew signal output
rlabel metal2 s 58254 0 58310 800 6 clk
port 3 nsew signal input
rlabel metal2 s 81622 0 81678 800 6 clk_en
port 4 nsew signal output
rlabel metal3 s 0 69912 800 70032 6 cs_en
port 5 nsew signal output
rlabel metal3 s 139200 23264 140000 23384 6 loopthrough_sel
port 6 nsew signal input
rlabel metal2 s 104898 139200 104954 140000 6 lt_sel_en
port 7 nsew signal output
rlabel metal3 s 139200 69912 140000 70032 6 minion_parity
port 8 nsew signal output
rlabel metal3 s 0 116560 800 116680 6 miso_en
port 9 nsew signal output
rlabel metal2 s 104898 0 104954 800 6 mosi_en
port 10 nsew signal output
rlabel metal2 s 128266 139200 128322 140000 6 mp_en
port 11 nsew signal output
rlabel metal2 s 11610 0 11666 800 6 reset
port 12 nsew signal input
rlabel metal2 s 34886 0 34942 800 6 reset_en
port 13 nsew signal output
rlabel metal2 s 128266 0 128322 800 6 sclk_en
port 14 nsew signal output
rlabel metal2 s 81622 139200 81678 140000 6 spi_min_cs
port 15 nsew signal input
rlabel metal2 s 34886 139200 34942 140000 6 spi_min_miso
port 16 nsew signal output
rlabel metal2 s 11610 139200 11666 140000 6 spi_min_mosi
port 17 nsew signal input
rlabel metal2 s 58254 139200 58310 140000 6 spi_min_sclk
port 18 nsew signal input
rlabel metal4 s 4208 2128 4528 137680 6 vccd1
port 19 nsew power input
rlabel metal4 s 34928 2128 35248 137680 6 vccd1
port 19 nsew power input
rlabel metal4 s 65648 2128 65968 137680 6 vccd1
port 19 nsew power input
rlabel metal4 s 96368 2128 96688 137680 6 vccd1
port 19 nsew power input
rlabel metal4 s 127088 2128 127408 137680 6 vccd1
port 19 nsew power input
rlabel metal4 s 19568 2128 19888 137680 6 vssd1
port 20 nsew ground input
rlabel metal4 s 50288 2128 50608 137680 6 vssd1
port 20 nsew ground input
rlabel metal4 s 81008 2128 81328 137680 6 vssd1
port 20 nsew ground input
rlabel metal4 s 111728 2128 112048 137680 6 vssd1
port 20 nsew ground input
<< properties >>
string FIXED_BBOX 0 0 140000 140000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 12025126
string GDS_FILE /home/acm289/ece5745-tapeout/openlane/project-group99/runs/project-group99/results/finishing/grp_99_SPI_TapeOutBlockRTL_32bits_5entries.magic.gds
string GDS_START 643446
<< end >>


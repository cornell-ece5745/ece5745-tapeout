magic
tech sky130A
magscale 1 2
timestamp 1655308115
<< obsli1 >>
rect 1104 2159 198812 197489
<< obsm1 >>
rect 14 2128 199718 197520
<< metal2 >>
rect 27066 199200 27122 200000
rect 70214 199200 70270 200000
rect 113362 199200 113418 200000
rect 156510 199200 156566 200000
rect 199658 199200 199714 200000
rect 18 0 74 800
rect 43166 0 43222 800
rect 86314 0 86370 800
rect 129462 0 129518 800
rect 172610 0 172666 800
<< obsm2 >>
rect 20 199144 27010 199322
rect 27178 199144 70158 199322
rect 70326 199144 113306 199322
rect 113474 199144 156454 199322
rect 156622 199144 199602 199322
rect 20 856 199712 199144
rect 130 800 43110 856
rect 43278 800 86258 856
rect 86426 800 129406 856
rect 129574 800 172554 856
rect 172722 800 199712 856
<< metal3 >>
rect 0 182248 800 182368
rect 199200 153688 200000 153808
rect 0 136688 800 136808
rect 199200 108128 200000 108248
rect 0 91128 800 91248
rect 199200 62568 200000 62688
rect 0 45568 800 45688
rect 199200 17008 200000 17128
<< obsm3 >>
rect 800 182448 199200 197505
rect 880 182168 199200 182448
rect 800 153888 199200 182168
rect 800 153608 199120 153888
rect 800 136888 199200 153608
rect 880 136608 199200 136888
rect 800 108328 199200 136608
rect 800 108048 199120 108328
rect 800 91328 199200 108048
rect 880 91048 199200 91328
rect 800 62768 199200 91048
rect 800 62488 199120 62768
rect 800 45768 199200 62488
rect 880 45488 199200 45768
rect 800 17208 199200 45488
rect 800 16928 199120 17208
rect 800 2143 199200 16928
<< metal4 >>
rect 4208 2128 4528 197520
rect 19568 2128 19888 197520
rect 34928 2128 35248 197520
rect 50288 2128 50608 197520
rect 65648 2128 65968 197520
rect 81008 2128 81328 197520
rect 96368 2128 96688 197520
rect 111728 2128 112048 197520
rect 127088 2128 127408 197520
rect 142448 2128 142768 197520
rect 157808 2128 158128 197520
rect 173168 2128 173488 197520
rect 188528 2128 188848 197520
<< obsm4 >>
rect 80651 76467 80928 143853
rect 81408 76467 96288 143853
rect 96768 76467 111648 143853
rect 112128 76467 127008 143853
rect 127488 76467 142368 143853
rect 142848 76467 154133 143853
<< labels >>
rlabel metal3 s 199200 17008 200000 17128 6 adapter_parity
port 1 nsew signal output
rlabel metal3 s 199200 153688 200000 153808 6 ap_en
port 2 nsew signal output
rlabel metal2 s 113362 199200 113418 200000 6 clk
port 3 nsew signal input
rlabel metal2 s 129462 0 129518 800 6 clk_en
port 4 nsew signal output
rlabel metal3 s 0 182248 800 182368 6 cs_en
port 5 nsew signal output
rlabel metal2 s 70214 199200 70270 200000 6 loopthrough_sel
port 6 nsew signal input
rlabel metal2 s 18 0 74 800 6 lt_sel_en
port 7 nsew signal output
rlabel metal2 s 199658 199200 199714 200000 6 minion_parity
port 8 nsew signal output
rlabel metal2 s 172610 0 172666 800 6 miso_en
port 9 nsew signal output
rlabel metal2 s 43166 0 43222 800 6 mosi_en
port 10 nsew signal output
rlabel metal3 s 0 45568 800 45688 6 mp_en
port 11 nsew signal output
rlabel metal3 s 199200 108128 200000 108248 6 reset
port 12 nsew signal input
rlabel metal3 s 0 91128 800 91248 6 reset_en
port 13 nsew signal output
rlabel metal2 s 156510 199200 156566 200000 6 sclk_en
port 14 nsew signal output
rlabel metal2 s 86314 0 86370 800 6 spi_min_cs
port 15 nsew signal input
rlabel metal3 s 0 136688 800 136808 6 spi_min_miso
port 16 nsew signal output
rlabel metal2 s 27066 199200 27122 200000 6 spi_min_mosi
port 17 nsew signal input
rlabel metal3 s 199200 62568 200000 62688 6 spi_min_sclk
port 18 nsew signal input
rlabel metal4 s 4208 2128 4528 197520 6 vccd1
port 19 nsew power input
rlabel metal4 s 34928 2128 35248 197520 6 vccd1
port 19 nsew power input
rlabel metal4 s 65648 2128 65968 197520 6 vccd1
port 19 nsew power input
rlabel metal4 s 96368 2128 96688 197520 6 vccd1
port 19 nsew power input
rlabel metal4 s 127088 2128 127408 197520 6 vccd1
port 19 nsew power input
rlabel metal4 s 157808 2128 158128 197520 6 vccd1
port 19 nsew power input
rlabel metal4 s 188528 2128 188848 197520 6 vccd1
port 19 nsew power input
rlabel metal4 s 19568 2128 19888 197520 6 vssd1
port 20 nsew ground input
rlabel metal4 s 50288 2128 50608 197520 6 vssd1
port 20 nsew ground input
rlabel metal4 s 81008 2128 81328 197520 6 vssd1
port 20 nsew ground input
rlabel metal4 s 111728 2128 112048 197520 6 vssd1
port 20 nsew ground input
rlabel metal4 s 142448 2128 142768 197520 6 vssd1
port 20 nsew ground input
rlabel metal4 s 173168 2128 173488 197520 6 vssd1
port 20 nsew ground input
<< properties >>
string FIXED_BBOX 0 0 200000 200000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 21142444
string GDS_FILE /home/acm289/ece5745-tapeout/openlane/project-group15/runs/project-group15/results/finishing/grp_15_SPI_TapeOutBlockRTL_32bits_5entries.magic.gds
string GDS_START 646196
<< end >>

